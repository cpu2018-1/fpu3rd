module fsqrt(
    input wire [31:0] x,
    output wire [31:0] y);

    function [36:0] TDATA (
	input [8:0] KEY
    );
    begin
        case(KEY)
        9'd256: TDATA = 37'b0000000000111111111100101111111111000;
        9'd257: TDATA = 37'b0000000010111111101100101111111101000;
        9'd258: TDATA = 37'b0000000100111111001100101111111011000;
        9'd259: TDATA = 37'b0000000110111110011101001111111001001;
        9'd260: TDATA = 37'b0000001000111101011110001111110111001;
        9'd261: TDATA = 37'b0000001010111100001111001111110101001;
        9'd262: TDATA = 37'b0000001100111010110000101111110011010;
        9'd263: TDATA = 37'b0000001110111001000011001111110001011;
        9'd264: TDATA = 37'b0000010000110111000110001111101111011;
        9'd265: TDATA = 37'b0000010010110100111001101111101101100;
        9'd266: TDATA = 37'b0000010100110010011110001111101011101;
        9'd267: TDATA = 37'b0000010110101111110011101111101001110;
        9'd268: TDATA = 37'b0000011000101100111010001111100111111;
        9'd269: TDATA = 37'b0000011010101001110001101111100110000;
        9'd270: TDATA = 37'b0000011100100110011010101111100100001;
        9'd271: TDATA = 37'b0000011110100010110100101111100010011;
        9'd272: TDATA = 37'b0000100000011111000000001111100000100;
        9'd273: TDATA = 37'b0000100010011010111101001111011110110;
        9'd274: TDATA = 37'b0000100100010110101011001111011100111;
        9'd275: TDATA = 37'b0000100110010010001011001111011011001;
        9'd276: TDATA = 37'b0000101000001101011100101111011001010;
        9'd277: TDATA = 37'b0000101010001000100000001111010111100;
        9'd278: TDATA = 37'b0000101100000011010101101111010101110;
        9'd279: TDATA = 37'b0000101101111101111100101111010100000;
        9'd280: TDATA = 37'b0000101111111000010101101111010010010;
        9'd281: TDATA = 37'b0000110001110010100000101111010000100;
        9'd282: TDATA = 37'b0000110011101100011101101111001110110;
        9'd283: TDATA = 37'b0000110101100110001101001111001101001;
        9'd284: TDATA = 37'b0000110111011111101111001111001011011;
        9'd285: TDATA = 37'b0000111001011001000011001111001001101;
        9'd286: TDATA = 37'b0000111011010010001001101111001000000;
        9'd287: TDATA = 37'b0000111101001011000010101111000110010;
        9'd288: TDATA = 37'b0000111111000011101110001111000100101;
        9'd289: TDATA = 37'b0001000000111100001100001111000010111;
        9'd290: TDATA = 37'b0001000010110100011100101111000001010;
        9'd291: TDATA = 37'b0001000100101100100000101110111111101;
        9'd292: TDATA = 37'b0001000110100100010110101110111110000;
        9'd293: TDATA = 37'b0001001000011100000000001110111100011;
        9'd294: TDATA = 37'b0001001010010011011100101110111010110;
        9'd295: TDATA = 37'b0001001100001010101011101110111001001;
        9'd296: TDATA = 37'b0001001110000001101110001110110111100;
        9'd297: TDATA = 37'b0001001111111000100011101110110101111;
        9'd298: TDATA = 37'b0001010001101111001100101110110100010;
        9'd299: TDATA = 37'b0001010011100101101000101110110010110;
        9'd300: TDATA = 37'b0001010101011011111000001110110001001;
        9'd301: TDATA = 37'b0001010111010001111011001110101111101;
        9'd302: TDATA = 37'b0001011001000111110001001110101110000;
        9'd303: TDATA = 37'b0001011010111101011011001110101100100;
        9'd304: TDATA = 37'b0001011100110010111000101110101010111;
        9'd305: TDATA = 37'b0001011110101000001001101110101001011;
        9'd306: TDATA = 37'b0001100000011101001110101110100111111;
        9'd307: TDATA = 37'b0001100010010010000111101110100110011;
        9'd308: TDATA = 37'b0001100100000110110100001110100100110;
        9'd309: TDATA = 37'b0001100101111011010100001110100011010;
        9'd310: TDATA = 37'b0001100111101111101000101110100001110;
        9'd311: TDATA = 37'b0001101001100011110001001110100000010;
        9'd312: TDATA = 37'b0001101011010111101101101110011110111;
        9'd313: TDATA = 37'b0001101101001011011110001110011101011;
        9'd314: TDATA = 37'b0001101110111111000011001110011011111;
        9'd315: TDATA = 37'b0001110000110010011100001110011010011;
        9'd316: TDATA = 37'b0001110010100101101001101110011001000;
        9'd317: TDATA = 37'b0001110100011000101011001110010111100;
        9'd318: TDATA = 37'b0001110110001011100001101110010110000;
        9'd319: TDATA = 37'b0001110111111110001100001110010100101;
        9'd320: TDATA = 37'b0001111001110000101011001110010011001;
        9'd321: TDATA = 37'b0001111011100010111111001110010001110;
        9'd322: TDATA = 37'b0001111101010101000111001110010000011;
        9'd323: TDATA = 37'b0001111111000111000100001110001110111;
        9'd324: TDATA = 37'b0010000000111000110110001110001101100;
        9'd325: TDATA = 37'b0010000010101010011100101110001100001;
        9'd326: TDATA = 37'b0010000100011011111000001110001010110;
        9'd327: TDATA = 37'b0010000110001101001000101110001001011;
        9'd328: TDATA = 37'b0010000111111110001101101110001000000;
        9'd329: TDATA = 37'b0010001001101111000111101110000110101;
        9'd330: TDATA = 37'b0010001011011111110111001110000101010;
        9'd331: TDATA = 37'b0010001101010000011011101110000011111;
        9'd332: TDATA = 37'b0010001111000000110101001110000010100;
        9'd333: TDATA = 37'b0010010000110001000011101110000001001;
        9'd334: TDATA = 37'b0010010010100001000111101101111111111;
        9'd335: TDATA = 37'b0010010100010001000001001101111110100;
        9'd336: TDATA = 37'b0010010110000000101111101101111101001;
        9'd337: TDATA = 37'b0010010111110000010011101101111011111;
        9'd338: TDATA = 37'b0010011001011111101100101101111010100;
        9'd339: TDATA = 37'b0010011011001110111011101101111001010;
        9'd340: TDATA = 37'b0010011100111110000000001101110111111;
        9'd341: TDATA = 37'b0010011110101100111010001101110110101;
        9'd342: TDATA = 37'b0010100000011011101001101101110101010;
        9'd343: TDATA = 37'b0010100010001010001110101101110100000;
        9'd344: TDATA = 37'b0010100011111000101001101101110010110;
        9'd345: TDATA = 37'b0010100101100110111010101101110001100;
        9'd346: TDATA = 37'b0010100111010101000000101101110000001;
        9'd347: TDATA = 37'b0010101001000010111101001101101110111;
        9'd348: TDATA = 37'b0010101010110000101111001101101101101;
        9'd349: TDATA = 37'b0010101100011110010111101101101100011;
        9'd350: TDATA = 37'b0010101110001011110101101101101011001;
        9'd351: TDATA = 37'b0010101111111001001001101101101001111;
        9'd352: TDATA = 37'b0010110001100110010011101101101000101;
        9'd353: TDATA = 37'b0010110011010011010100001101100111011;
        9'd354: TDATA = 37'b0010110101000000001010101101100110001;
        9'd355: TDATA = 37'b0010110110101100110111001101100101000;
        9'd356: TDATA = 37'b0010111000011001011010001101100011110;
        9'd357: TDATA = 37'b0010111010000101110011001101100010100;
        9'd358: TDATA = 37'b0010111011110010000010001101100001011;
        9'd359: TDATA = 37'b0010111101011110001000001101100000001;
        9'd360: TDATA = 37'b0010111111001010000100001101011110111;
        9'd361: TDATA = 37'b0011000000110101110110101101011101110;
        9'd362: TDATA = 37'b0011000010100001011111101101011100100;
        9'd363: TDATA = 37'b0011000100001100111111001101011011011;
        9'd364: TDATA = 37'b0011000101111000010101001101011010001;
        9'd365: TDATA = 37'b0011000111100011100001101101011001000;
        9'd366: TDATA = 37'b0011001001001110100101001101010111111;
        9'd367: TDATA = 37'b0011001010111001011111001101010110101;
        9'd368: TDATA = 37'b0011001100100100001111101101010101100;
        9'd369: TDATA = 37'b0011001110001110110111001101010100011;
        9'd370: TDATA = 37'b0011001111111001010101001101010011010;
        9'd371: TDATA = 37'b0011010001100011101010001101010010000;
        9'd372: TDATA = 37'b0011010011001101110101101101010000111;
        9'd373: TDATA = 37'b0011010100110111111000101101001111110;
        9'd374: TDATA = 37'b0011010110100001110010001101001110101;
        9'd375: TDATA = 37'b0011011000001011100010101101001101100;
        9'd376: TDATA = 37'b0011011001110101001010001101001100011;
        9'd377: TDATA = 37'b0011011011011110101000101101001011010;
        9'd378: TDATA = 37'b0011011101000111111110001101001010001;
        9'd379: TDATA = 37'b0011011110110001001011001101001001000;
        9'd380: TDATA = 37'b0011100000011010001110101101000111111;
        9'd381: TDATA = 37'b0011100010000011001001101101000110111;
        9'd382: TDATA = 37'b0011100011101011111100001101000101110;
        9'd383: TDATA = 37'b0011100101010100100101101101000100101;
        9'd384: TDATA = 37'b0011100110111101000110001101000011100;
        9'd385: TDATA = 37'b0011101000100101011110001101000010100;
        9'd386: TDATA = 37'b0011101010001101101101101101000001011;
        9'd387: TDATA = 37'b0011101011110101110100101101000000010;
        9'd388: TDATA = 37'b0011101101011101110010101100111111010;
        9'd389: TDATA = 37'b0011101111000101101000001100111110001;
        9'd390: TDATA = 37'b0011110000101101010101001100111101001;
        9'd391: TDATA = 37'b0011110010010100111010001100111100000;
        9'd392: TDATA = 37'b0011110011111100010110001100111011000;
        9'd393: TDATA = 37'b0011110101100011101001101100111010000;
        9'd394: TDATA = 37'b0011110111001010110101001100111000111;
        9'd395: TDATA = 37'b0011111000110001111000001100110111111;
        9'd396: TDATA = 37'b0011111010011000110010101100110110110;
        9'd397: TDATA = 37'b0011111011111111100101001100110101110;
        9'd398: TDATA = 37'b0011111101100110001111001100110100110;
        9'd399: TDATA = 37'b0011111111001100110000101100110011110;
        9'd400: TDATA = 37'b0100000000110011001010101100110010110;
        9'd401: TDATA = 37'b0100000010011001011011101100110001101;
        9'd402: TDATA = 37'b0100000011111111100101001100110000101;
        9'd403: TDATA = 37'b0100000101100101100110001100101111101;
        9'd404: TDATA = 37'b0100000111001011011111001100101110101;
        9'd405: TDATA = 37'b0100001000110001010000001100101101101;
        9'd406: TDATA = 37'b0100001010010110111001001100101100101;
        9'd407: TDATA = 37'b0100001011111100011010001100101011101;
        9'd408: TDATA = 37'b0100001101100001110011101100101010101;
        9'd409: TDATA = 37'b0100001111000111000100101100101001101;
        9'd410: TDATA = 37'b0100010000101100001101101100101000101;
        9'd411: TDATA = 37'b0100010010010001001111001100100111101;
        9'd412: TDATA = 37'b0100010011110110001000101100100110110;
        9'd413: TDATA = 37'b0100010101011010111010001100100101110;
        9'd414: TDATA = 37'b0100010110111111100100001100100100110;
        9'd415: TDATA = 37'b0100011000100100000110001100100011110;
        9'd416: TDATA = 37'b0100011010001000100000001100100010110;
        9'd417: TDATA = 37'b0100011011101100110011001100100001111;
        9'd418: TDATA = 37'b0100011101010000111110001100100000111;
        9'd419: TDATA = 37'b0100011110110101000001001100011111111;
        9'd420: TDATA = 37'b0100100000011000111100101100011111000;
        9'd421: TDATA = 37'b0100100001111100110001001100011110000;
        9'd422: TDATA = 37'b0100100011100000011101001100011101001;
        9'd423: TDATA = 37'b0100100101000100000010001100011100001;
        9'd424: TDATA = 37'b0100100110100111011111101100011011010;
        9'd425: TDATA = 37'b0100101000001010110101101100011010010;
        9'd426: TDATA = 37'b0100101001101110000100001100011001011;
        9'd427: TDATA = 37'b0100101011010001001011001100011000011;
        9'd428: TDATA = 37'b0100101100110100001010101100010111100;
        9'd429: TDATA = 37'b0100101110010111000011001100010110101;
        9'd430: TDATA = 37'b0100101111111001110011101100010101101;
        9'd431: TDATA = 37'b0100110001011100011101001100010100110;
        9'd432: TDATA = 37'b0100110010111110111111101100010011111;
        9'd433: TDATA = 37'b0100110100100001011010101100010010111;
        9'd434: TDATA = 37'b0100110110000011101110001100010010000;
        9'd435: TDATA = 37'b0100110111100101111010101100010001001;
        9'd436: TDATA = 37'b0100111001000111111111101100010000010;
        9'd437: TDATA = 37'b0100111010101001111101101100001111010;
        9'd438: TDATA = 37'b0100111100001011110100101100001110011;
        9'd439: TDATA = 37'b0100111101101101100100001100001101100;
        9'd440: TDATA = 37'b0100111111001111001101001100001100101;
        9'd441: TDATA = 37'b0101000000110000101110101100001011110;
        9'd442: TDATA = 37'b0101000010010010001001001100001010111;
        9'd443: TDATA = 37'b0101000011110011011100101100001010000;
        9'd444: TDATA = 37'b0101000101010100101000101100001001001;
        9'd445: TDATA = 37'b0101000110110101101110001100001000010;
        9'd446: TDATA = 37'b0101001000010110101100101100000111011;
        9'd447: TDATA = 37'b0101001001110111100100001100000110100;
        9'd448: TDATA = 37'b0101001011011000010100101100000101101;
        9'd449: TDATA = 37'b0101001100111000111110001100000100110;
        9'd450: TDATA = 37'b0101001110011001100001001100000011111;
        9'd451: TDATA = 37'b0101001111111001111101001100000011001;
        9'd452: TDATA = 37'b0101010001011010010010001100000010010;
        9'd453: TDATA = 37'b0101010010111010100000101100000001011;
        9'd454: TDATA = 37'b0101010100011010101000001100000000100;
        9'd455: TDATA = 37'b0101010101111010101000101011111111101;
        9'd456: TDATA = 37'b0101010111011010100010101011111110111;
        9'd457: TDATA = 37'b0101011000111010010110001011111110000;
        9'd458: TDATA = 37'b0101011010011010000010101011111101001;
        9'd459: TDATA = 37'b0101011011111001101000101011111100011;
        9'd460: TDATA = 37'b0101011101011001000111101011111011100;
        9'd461: TDATA = 37'b0101011110111000100000101011111010101;
        9'd462: TDATA = 37'b0101100000010111110010101011111001111;
        9'd463: TDATA = 37'b0101100001110110111110001011111001000;
        9'd464: TDATA = 37'b0101100011010110000010101011111000010;
        9'd465: TDATA = 37'b0101100100110101000001001011110111011;
        9'd466: TDATA = 37'b0101100110010011111001001011110110101;
        9'd467: TDATA = 37'b0101100111110010101010001011110101110;
        9'd468: TDATA = 37'b0101101001010001010101001011110101000;
        9'd469: TDATA = 37'b0101101010101111111001001011110100001;
        9'd470: TDATA = 37'b0101101100001110010111001011110011011;
        9'd471: TDATA = 37'b0101101101101100101110101011110010100;
        9'd472: TDATA = 37'b0101101111001010111111101011110001110;
        9'd473: TDATA = 37'b0101110000101001001010101011110001000;
        9'd474: TDATA = 37'b0101110010000111001110101011110000001;
        9'd475: TDATA = 37'b0101110011100101001100101011101111011;
        9'd476: TDATA = 37'b0101110101000011000100101011101110101;
        9'd477: TDATA = 37'b0101110110100000110110001011101101110;
        9'd478: TDATA = 37'b0101110111111110100001001011101101000;
        9'd479: TDATA = 37'b0101111001011100000101101011101100010;
        9'd480: TDATA = 37'b0101111010111001100100101011101011011;
        9'd481: TDATA = 37'b0101111100010110111100101011101010101;
        9'd482: TDATA = 37'b0101111101110100001111001011101001111;
        9'd483: TDATA = 37'b0101111111010001011011001011101001001;
        9'd484: TDATA = 37'b0110000000101110100000101011101000011;
        9'd485: TDATA = 37'b0110000010001011100000101011100111101;
        9'd486: TDATA = 37'b0110000011101000011010001011100110110;
        9'd487: TDATA = 37'b0110000101000101001101101011100110000;
        9'd488: TDATA = 37'b0110000110100001111010101011100101010;
        9'd489: TDATA = 37'b0110000111111110100010001011100100100;
        9'd490: TDATA = 37'b0110001001011011000011001011100011110;
        9'd491: TDATA = 37'b0110001010110111011110101011100011000;
        9'd492: TDATA = 37'b0110001100010011110011101011100010010;
        9'd493: TDATA = 37'b0110001101110000000010101011100001100;
        9'd494: TDATA = 37'b0110001111001100001100001011100000110;
        9'd495: TDATA = 37'b0110010000101000001111001011100000000;
        9'd496: TDATA = 37'b0110010010000100001100101011011111010;
        9'd497: TDATA = 37'b0110010011100000000100001011011110100;
        9'd498: TDATA = 37'b0110010100111011110101101011011101111;
        9'd499: TDATA = 37'b0110010110010111100001001011011101001;
        9'd500: TDATA = 37'b0110010111110011000110101011011100011;
        9'd501: TDATA = 37'b0110011001001110100110101011011011101;
        9'd502: TDATA = 37'b0110011010101010000000101011011010111;
        9'd503: TDATA = 37'b0110011100000101010101001011011010001;
        9'd504: TDATA = 37'b0110011101100000100011001011011001100;
        9'd505: TDATA = 37'b0110011110111011101100001011011000110;
        9'd506: TDATA = 37'b0110100000010110101110101011011000000;
        9'd507: TDATA = 37'b0110100001110001101100001011010111010;
        9'd508: TDATA = 37'b0110100011001100100011001011010110101;
        9'd509: TDATA = 37'b0110100100100111010101001011010101111;
        9'd510: TDATA = 37'b0110100110000010000001001011010101001;
        9'd511: TDATA = 37'b0110100111011100100111001011010100011;
        9'd0: TDATA = 37'b0110101001100100010110010110100110110;
        9'd1: TDATA = 37'b0110101100011001000000110110100011111;
        9'd2: TDATA = 37'b0110101111001101010101010110100001001;
        9'd3: TDATA = 37'b0110110010000001010011010110011110011;
        9'd4: TDATA = 37'b0110110100110100111010110110011011101;
        9'd5: TDATA = 37'b0110110111101000001100110110011000111;
        9'd6: TDATA = 37'b0110111010011011001000010110010110001;
        9'd7: TDATA = 37'b0110111101001101101110010110010011011;
        9'd8: TDATA = 37'b0110111111111111111110110110010000110;
        9'd9: TDATA = 37'b0111000010110001111001110110001110000;
        9'd10: TDATA = 37'b0111000101100011011110110110001011011;
        9'd11: TDATA = 37'b0111001000010100101111010110001000101;
        9'd12: TDATA = 37'b0111001011000101101001110110000110000;
        9'd13: TDATA = 37'b0111001101110110001111110110000011011;
        9'd14: TDATA = 37'b0111010000100110100000110110000000110;
        9'd15: TDATA = 37'b0111010011010110011100110101111110010;
        9'd16: TDATA = 37'b0111010110000110000100010101111011101;
        9'd17: TDATA = 37'b0111011000110101010110110101111001000;
        9'd18: TDATA = 37'b0111011011100100010101010101110110100;
        9'd19: TDATA = 37'b0111011110010010111110110101110100000;
        9'd20: TDATA = 37'b0111100001000001010100010101110001011;
        9'd21: TDATA = 37'b0111100011101111010101110101101110111;
        9'd22: TDATA = 37'b0111100110011101000011010101101100011;
        9'd23: TDATA = 37'b0111101001001010011100110101101010000;
        9'd24: TDATA = 37'b0111101011110111100010010101100111100;
        9'd25: TDATA = 37'b0111101110100100010100010101100101000;
        9'd26: TDATA = 37'b0111110001010000110010010101100010100;
        9'd27: TDATA = 37'b0111110011111100111101010101100000001;
        9'd28: TDATA = 37'b0111110110101000110100110101011101110;
        9'd29: TDATA = 37'b0111111001010100011000110101011011010;
        9'd30: TDATA = 37'b0111111011111111101001010101011000111;
        9'd31: TDATA = 37'b0111111110101010100111010101010110100;
        9'd32: TDATA = 37'b1000000001010101010001110101010100001;
        9'd33: TDATA = 37'b1000000011111111101001010101010001110;
        9'd34: TDATA = 37'b1000000110101001101110010101001111100;
        9'd35: TDATA = 37'b1000001001010011100000110101001101001;
        9'd36: TDATA = 37'b1000001011111101000000010101001010110;
        9'd37: TDATA = 37'b1000001110100110001101010101001000100;
        9'd38: TDATA = 37'b1000010001001111000111110101000110001;
        9'd39: TDATA = 37'b1000010011110111110000010101000011111;
        9'd40: TDATA = 37'b1000010110100000000110010101000001101;
        9'd41: TDATA = 37'b1000011001001000001010010100111111011;
        9'd42: TDATA = 37'b1000011011101111111100010100111101001;
        9'd43: TDATA = 37'b1000011110010111011011110100111010111;
        9'd44: TDATA = 37'b1000100000111110101001110100111000101;
        9'd45: TDATA = 37'b1000100011100101100110010100110110011;
        9'd46: TDATA = 37'b1000100110001100010000110100110100010;
        9'd47: TDATA = 37'b1000101000110010101001010100110010000;
        9'd48: TDATA = 37'b1000101011011000110000110100101111111;
        9'd49: TDATA = 37'b1000101101111110100110110100101101101;
        9'd50: TDATA = 37'b1000110000100100001011010100101011100;
        9'd51: TDATA = 37'b1000110011001001011110110100101001011;
        9'd52: TDATA = 37'b1000110101101110100000110100100111010;
        9'd53: TDATA = 37'b1000111000010011010001110100100101000;
        9'd54: TDATA = 37'b1000111010110111110001110100100010111;
        9'd55: TDATA = 37'b1000111101011100000000110100100000111;
        9'd56: TDATA = 37'b1000111111111111111110110100011110110;
        9'd57: TDATA = 37'b1001000010100011101100010100011100101;
        9'd58: TDATA = 37'b1001000101000111001000110100011010100;
        9'd59: TDATA = 37'b1001000111101010010100110100011000100;
        9'd60: TDATA = 37'b1001001010001101010000010100010110011;
        9'd61: TDATA = 37'b1001001100101111111011010100010100011;
        9'd62: TDATA = 37'b1001001111010010010110010100010010011;
        9'd63: TDATA = 37'b1001010001110100100000110100010000010;
        9'd64: TDATA = 37'b1001010100010110011010110100001110010;
        9'd65: TDATA = 37'b1001010110111000000100110100001100010;
        9'd66: TDATA = 37'b1001011001011001011110110100001010010;
        9'd67: TDATA = 37'b1001011011111010101000110100001000010;
        9'd68: TDATA = 37'b1001011110011011100010110100000110010;
        9'd69: TDATA = 37'b1001100000111100001100110100000100010;
        9'd70: TDATA = 37'b1001100011011100100111010100000010010;
        9'd71: TDATA = 37'b1001100101111100110001110100000000011;
        9'd72: TDATA = 37'b1001101000011100101100110011111110011;
        9'd73: TDATA = 37'b1001101010111100011000010011111100100;
        9'd74: TDATA = 37'b1001101101011011110100010011111010100;
        9'd75: TDATA = 37'b1001101111111011000000110011111000101;
        9'd76: TDATA = 37'b1001110010011001111101110011110110110;
        9'd77: TDATA = 37'b1001110100111000101011110011110100110;
        9'd78: TDATA = 37'b1001110111010111001010010011110010111;
        9'd79: TDATA = 37'b1001111001110101011001110011110001000;
        9'd80: TDATA = 37'b1001111100010011011010010011101111001;
        9'd81: TDATA = 37'b1001111110110001001011110011101101010;
        9'd82: TDATA = 37'b1010000001001110101110010011101011011;
        9'd83: TDATA = 37'b1010000011101100000001110011101001100;
        9'd84: TDATA = 37'b1010000110001001000110010011100111101;
        9'd85: TDATA = 37'b1010001000100101111100010011100101111;
        9'd86: TDATA = 37'b1010001011000010100011110011100100000;
        9'd87: TDATA = 37'b1010001101011110111100110011100010001;
        9'd88: TDATA = 37'b1010001111111011000110110011100000011;
        9'd89: TDATA = 37'b1010010010010111000010010011011110100;
        9'd90: TDATA = 37'b1010010100110010101111110011011100110;
        9'd91: TDATA = 37'b1010010111001110001110010011011011000;
        9'd92: TDATA = 37'b1010011001101001011110110011011001001;
        9'd93: TDATA = 37'b1010011100000100100001010011010111011;
        9'd94: TDATA = 37'b1010011110011111010101010011010101101;
        9'd95: TDATA = 37'b1010100000111001111011010011010011111;
        9'd96: TDATA = 37'b1010100011010100010011010011010010001;
        9'd97: TDATA = 37'b1010100101101110011101010011010000011;
        9'd98: TDATA = 37'b1010101000001000011001010011001110101;
        9'd99: TDATA = 37'b1010101010100010000111010011001100111;
        9'd100: TDATA = 37'b1010101100111011100111110011001011001;
        9'd101: TDATA = 37'b1010101111010100111010010011001001100;
        9'd102: TDATA = 37'b1010110001101101111110110011000111110;
        9'd103: TDATA = 37'b1010110100000110110101110011000110000;
        9'd104: TDATA = 37'b1010110110011111011111010011000100011;
        9'd105: TDATA = 37'b1010111000110111111011010011000010101;
        9'd106: TDATA = 37'b1010111011010000001001110011000001000;
        9'd107: TDATA = 37'b1010111101101000001011010010111111010;
        9'd108: TDATA = 37'b1010111111111111111110110010111101101;
        9'd109: TDATA = 37'b1011000010010111100101010010111100000;
        9'd110: TDATA = 37'b1011000100101110111110010010111010011;
        9'd111: TDATA = 37'b1011000111000110001010010010111000101;
        9'd112: TDATA = 37'b1011001001011101001000110010110111000;
        9'd113: TDATA = 37'b1011001011110011111010110010110101011;
        9'd114: TDATA = 37'b1011001110001010011111010010110011110;
        9'd115: TDATA = 37'b1011010000100000110110110010110010001;
        9'd116: TDATA = 37'b1011010010110111000001010010110000100;
        9'd117: TDATA = 37'b1011010101001100111111010010101110111;
        9'd118: TDATA = 37'b1011010111100010110000010010101101011;
        9'd119: TDATA = 37'b1011011001111000010100010010101011110;
        9'd120: TDATA = 37'b1011011100001101101011110010101010001;
        9'd121: TDATA = 37'b1011011110100010110110010010101000100;
        9'd122: TDATA = 37'b1011100000110111110100110010100111000;
        9'd123: TDATA = 37'b1011100011001100100110010010100101011;
        9'd124: TDATA = 37'b1011100101100001001011010010100011111;
        9'd125: TDATA = 37'b1011100111110101100011010010100010010;
        9'd126: TDATA = 37'b1011101010001001101111110010100000110;
        9'd127: TDATA = 37'b1011101100011101101111010010011111001;
        9'd128: TDATA = 37'b1011101110110001100010010010011101101;
        9'd129: TDATA = 37'b1011110001000101001001110010011100001;
        9'd130: TDATA = 37'b1011110011011000100100010010011010101;
        9'd131: TDATA = 37'b1011110101101011110010110010011001000;
        9'd132: TDATA = 37'b1011110111111110110101010010010111100;
        9'd133: TDATA = 37'b1011111010010001101011110010010110000;
        9'd134: TDATA = 37'b1011111100100100010101110010010100100;
        9'd135: TDATA = 37'b1011111110110110110100010010010011000;
        9'd136: TDATA = 37'b1100000001001001000110010010010001100;
        9'd137: TDATA = 37'b1100000011011011001100110010010000000;
        9'd138: TDATA = 37'b1100000101101101000111010010001110101;
        9'd139: TDATA = 37'b1100000111111110110101110010001101001;
        9'd140: TDATA = 37'b1100001010010000011000110010001011101;
        9'd141: TDATA = 37'b1100001100100001101111110010001010001;
        9'd142: TDATA = 37'b1100001110110010111011010010001000110;
        9'd143: TDATA = 37'b1100010001000011111011010010000111010;
        9'd144: TDATA = 37'b1100010011010100101111010010000101110;
        9'd145: TDATA = 37'b1100010101100101011000010010000100011;
        9'd146: TDATA = 37'b1100010111110101110101010010000010111;
        9'd147: TDATA = 37'b1100011010000110000110110010000001100;
        9'd148: TDATA = 37'b1100011100010110001100110010000000000;
        9'd149: TDATA = 37'b1100011110100110000111110001111110101;
        9'd150: TDATA = 37'b1100100000110101110111010001111101010;
        9'd151: TDATA = 37'b1100100011000101011011010001111011111;
        9'd152: TDATA = 37'b1100100101010100110100010001111010011;
        9'd153: TDATA = 37'b1100100111100100000001110001111001000;
        9'd154: TDATA = 37'b1100101001110011000100010001110111101;
        9'd155: TDATA = 37'b1100101100000001111011110001110110010;
        9'd156: TDATA = 37'b1100101110010000100111110001110100111;
        9'd157: TDATA = 37'b1100110000011111001001010001110011100;
        9'd158: TDATA = 37'b1100110010101101011111010001110010001;
        9'd159: TDATA = 37'b1100110100111011101010010001110000110;
        9'd160: TDATA = 37'b1100110111001001101010110001101111011;
        9'd161: TDATA = 37'b1100111001010111011111110001101110000;
        9'd162: TDATA = 37'b1100111011100101001010010001101100101;
        9'd163: TDATA = 37'b1100111101110010101001110001101011010;
        9'd164: TDATA = 37'b1100111111111111111110110001101001111;
        9'd165: TDATA = 37'b1101000010001101001000110001101000101;
        9'd166: TDATA = 37'b1101000100011010001000010001100111010;
        9'd167: TDATA = 37'b1101000110100110111100110001100101111;
        9'd168: TDATA = 37'b1101001000110011100110110001100100101;
        9'd169: TDATA = 37'b1101001011000000000110010001100011010;
        9'd170: TDATA = 37'b1101001101001100011011010001100010000;
        9'd171: TDATA = 37'b1101001111011000100101110001100000101;
        9'd172: TDATA = 37'b1101010001100100100101110001011111011;
        9'd173: TDATA = 37'b1101010011110000011011010001011110000;
        9'd174: TDATA = 37'b1101010101111100000110010001011100110;
        9'd175: TDATA = 37'b1101011000000111100110110001011011011;
        9'd176: TDATA = 37'b1101011010010010111101010001011010001;
        9'd177: TDATA = 37'b1101011100011110001001010001011000111;
        9'd178: TDATA = 37'b1101011110101001001010110001010111101;
        9'd179: TDATA = 37'b1101100000110100000010010001010110010;
        9'd180: TDATA = 37'b1101100010111110101111110001010101000;
        9'd181: TDATA = 37'b1101100101001001010010110001010011110;
        9'd182: TDATA = 37'b1101100111010011101011110001010010100;
        9'd183: TDATA = 37'b1101101001011101111010110001010001010;
        9'd184: TDATA = 37'b1101101011100111111111110001010000000;
        9'd185: TDATA = 37'b1101101101110001111010110001001110110;
        9'd186: TDATA = 37'b1101101111111011101011010001001101100;
        9'd187: TDATA = 37'b1101110010000101010010010001001100010;
        9'd188: TDATA = 37'b1101110100001110101111010001001011000;
        9'd189: TDATA = 37'b1101110110011000000010010001001001110;
        9'd190: TDATA = 37'b1101111000100001001011110001001000100;
        9'd191: TDATA = 37'b1101111010101010001010110001000111011;
        9'd192: TDATA = 37'b1101111100110011000000110001000110001;
        9'd193: TDATA = 37'b1101111110111011101100010001000100111;
        9'd194: TDATA = 37'b1110000001000100001110110001000011101;
        9'd195: TDATA = 37'b1110000011001100100111010001000010100;
        9'd196: TDATA = 37'b1110000101010100110101110001000001010;
        9'd197: TDATA = 37'b1110000111011100111010110001000000000;
        9'd198: TDATA = 37'b1110001001100100110110110000111110111;
        9'd199: TDATA = 37'b1110001011101100101000110000111101101;
        9'd200: TDATA = 37'b1110001101110100010000110000111100100;
        9'd201: TDATA = 37'b1110001111111011101111110000111011010;
        9'd202: TDATA = 37'b1110010010000011000101010000111010001;
        9'd203: TDATA = 37'b1110010100001010010001010000111000111;
        9'd204: TDATA = 37'b1110010110010001010100010000110111110;
        9'd205: TDATA = 37'b1110011000011000001101010000110110101;
        9'd206: TDATA = 37'b1110011010011110111101010000110101011;
        9'd207: TDATA = 37'b1110011100100101100011110000110100010;
        9'd208: TDATA = 37'b1110011110101100000001010000110011001;
        9'd209: TDATA = 37'b1110100000110010010101010000110001111;
        9'd210: TDATA = 37'b1110100010111000011111110000110000110;
        9'd211: TDATA = 37'b1110100100111110100001110000101111101;
        9'd212: TDATA = 37'b1110100111000100011010010000101110100;
        9'd213: TDATA = 37'b1110101001001010001001010000101101011;
        9'd214: TDATA = 37'b1110101011001111101111110000101100010;
        9'd215: TDATA = 37'b1110101101010101001100110000101011001;
        9'd216: TDATA = 37'b1110101111011010100000110000101010000;
        9'd217: TDATA = 37'b1110110001011111101011110000101000111;
        9'd218: TDATA = 37'b1110110011100100101101110000100111110;
        9'd219: TDATA = 37'b1110110101101001100110110000100110101;
        9'd220: TDATA = 37'b1110110111101110010111010000100101100;
        9'd221: TDATA = 37'b1110111001110010111110010000100100011;
        9'd222: TDATA = 37'b1110111011110111011100110000100011010;
        9'd223: TDATA = 37'b1110111101111011110010010000100010001;
        9'd224: TDATA = 37'b1110111111111111111110110000100001000;
        9'd225: TDATA = 37'b1111000010000100000010110000011111111;
        9'd226: TDATA = 37'b1111000100000111111101110000011110111;
        9'd227: TDATA = 37'b1111000110001011110000010000011101110;
        9'd228: TDATA = 37'b1111001000001111011001110000011100101;
        9'd229: TDATA = 37'b1111001010010010111010110000011011101;
        9'd230: TDATA = 37'b1111001100010110010010110000011010100;
        9'd231: TDATA = 37'b1111001110011001100010110000011001011;
        9'd232: TDATA = 37'b1111010000011100101001110000011000011;
        9'd233: TDATA = 37'b1111010010011111100111110000010111010;
        9'd234: TDATA = 37'b1111010100100010011101110000010110010;
        9'd235: TDATA = 37'b1111010110100101001011010000010101001;
        9'd236: TDATA = 37'b1111011000100111110000010000010100001;
        9'd237: TDATA = 37'b1111011010101010001100010000010011000;
        9'd238: TDATA = 37'b1111011100101100100000010000010010000;
        9'd239: TDATA = 37'b1111011110101110101011110000010000111;
        9'd240: TDATA = 37'b1111100000110000101110110000001111111;
        9'd241: TDATA = 37'b1111100010110010101001110000001110111;
        9'd242: TDATA = 37'b1111100100110100011011110000001101110;
        9'd243: TDATA = 37'b1111100110110110000110010000001100110;
        9'd244: TDATA = 37'b1111101000110111100111110000001011110;
        9'd245: TDATA = 37'b1111101010111001000001010000001010101;
        9'd246: TDATA = 37'b1111101100111010010010010000001001101;
        9'd247: TDATA = 37'b1111101110111011011011010000001000101;
        9'd248: TDATA = 37'b1111110000111100011100010000000111101;
        9'd249: TDATA = 37'b1111110010111101010100110000000110101;
        9'd250: TDATA = 37'b1111110100111110000101010000000101100;
        9'd251: TDATA = 37'b1111110110111110101101010000000100100;
        9'd252: TDATA = 37'b1111111000111111001101110000000011100;
        9'd253: TDATA = 37'b1111111010111111100101110000000010100;
        9'd254: TDATA = 37'b1111111100111111110101110000000001100;
        9'd255: TDATA = 37'b1111111110111111111101110000000000100;
        endcase
    end
    endfunction

    wire [7:0] ex;
    assign ex = x[30:23];
    
    wire [8:0] key;
    wire pm;
    wire [13:0] h;
    assign key = x[23:15];
    assign pm = x[14];
    assign h = x[13:0];

    wire [36:0] tdata;
    assign tdata = TDATA(key);

    wire [22:0] rtx0;
    wire [13:0] rtx0_inv;
    assign rtx0 = tdata[36:14];
    assign rtx0_inv = tdata[13:0];

    wire check_zero;
    assign check_zero = (x[30:0] == 31'b0);

    wire [7:0] ey;
    assign ey = (check_zero) ? 8'b0: 8'd63 + ex[7:1] + ex[0];

    wire [13:0] noth;
    assign noth = ~h;

    wire [36:0] my_extend1;
    assign my_extend1 = {rtx0,14'b0} + rtx0_inv * h;

    wire [36:0] my_extend2;
    assign my_extend2 = {rtx0,14'b0} - rtx0_inv * noth;

    wire [22:0] my;
    assign my = (pm) ? my_extend1[36:14]: my_extend2[36:14];

    assign y = {1'b0,ey,my};

endmodule

