module fsqrt(
    input wire [31:0] x,
    output wire [31:0] y);

    function [36:0] TDATA (
	input [9:0] KEY
    );
    begin
        case(KEY)
        10'd512: TDATA = 37'b0000000000000000000000010000000000000;
        10'd513: TDATA = 37'b0000000000111111111110001111111111000;
        10'd514: TDATA = 37'b0000000001111111111000001111111110000;
        10'd515: TDATA = 37'b0000000010111111101110001111111101000;
        10'd516: TDATA = 37'b0000000011111111100000001111111100000;
        10'd517: TDATA = 37'b0000000100111111001110001111111011000;
        10'd518: TDATA = 37'b0000000101111110111000101111111010000;
        10'd519: TDATA = 37'b0000000110111110011110101111111001001;
        10'd520: TDATA = 37'b0000000111111110000001001111111000001;
        10'd521: TDATA = 37'b0000001000111101011111101111110111001;
        10'd522: TDATA = 37'b0000001001111100111010001111110110001;
        10'd523: TDATA = 37'b0000001010111100010000101111110101001;
        10'd524: TDATA = 37'b0000001011111011100011101111110100010;
        10'd525: TDATA = 37'b0000001100111010110010001111110011010;
        10'd526: TDATA = 37'b0000001101111001111101101111110010010;
        10'd527: TDATA = 37'b0000001110111001000100101111110001011;
        10'd528: TDATA = 37'b0000001111111000001000001111110000011;
        10'd529: TDATA = 37'b0000010000110111000111101111101111011;
        10'd530: TDATA = 37'b0000010001110110000011001111101110100;
        10'd531: TDATA = 37'b0000010010110100111011001111101101100;
        10'd532: TDATA = 37'b0000010011110011101111101111101100101;
        10'd533: TDATA = 37'b0000010100110010011111101111101011101;
        10'd534: TDATA = 37'b0000010101110001001100101111101010101;
        10'd535: TDATA = 37'b0000010110101111110101001111101001110;
        10'd536: TDATA = 37'b0000010111101110011010001111101000110;
        10'd537: TDATA = 37'b0000011000101100111011101111100111111;
        10'd538: TDATA = 37'b0000011001101011011001101111100111000;
        10'd539: TDATA = 37'b0000011010101001110011001111100110000;
        10'd540: TDATA = 37'b0000011011101000001001101111100101001;
        10'd541: TDATA = 37'b0000011100100110011100001111100100001;
        10'd542: TDATA = 37'b0000011101100100101011001111100011010;
        10'd543: TDATA = 37'b0000011110100010110110001111100010011;
        10'd544: TDATA = 37'b0000011111100000111101101111100001011;
        10'd545: TDATA = 37'b0000100000011111000001101111100000100;
        10'd546: TDATA = 37'b0000100001011101000001101111011111101;
        10'd547: TDATA = 37'b0000100010011010111110101111011110110;
        10'd548: TDATA = 37'b0000100011011000110111101111011101110;
        10'd549: TDATA = 37'b0000100100010110101100101111011100111;
        10'd550: TDATA = 37'b0000100101010100011110101111011100000;
        10'd551: TDATA = 37'b0000100110010010001100101111011011001;
        10'd552: TDATA = 37'b0000100111001111110111001111011010010;
        10'd553: TDATA = 37'b0000101000001101011110001111011001010;
        10'd554: TDATA = 37'b0000101001001011000001101111011000011;
        10'd555: TDATA = 37'b0000101010001000100001101111010111100;
        10'd556: TDATA = 37'b0000101011000101111110001111010110101;
        10'd557: TDATA = 37'b0000101100000011010111001111010101110;
        10'd558: TDATA = 37'b0000101101000000101100001111010100111;
        10'd559: TDATA = 37'b0000101101111101111110001111010100000;
        10'd560: TDATA = 37'b0000101110111011001100001111010011001;
        10'd561: TDATA = 37'b0000101111111000010111001111010010010;
        10'd562: TDATA = 37'b0000110000110101011110001111010001011;
        10'd563: TDATA = 37'b0000110001110010100010001111010000100;
        10'd564: TDATA = 37'b0000110010101111100010101111001111101;
        10'd565: TDATA = 37'b0000110011101100011111001111001110110;
        10'd566: TDATA = 37'b0000110100101001011000101111001101111;
        10'd567: TDATA = 37'b0000110101100110001110101111001101001;
        10'd568: TDATA = 37'b0000110110100011000001001111001100010;
        10'd569: TDATA = 37'b0000110111011111110000101111001011011;
        10'd570: TDATA = 37'b0000111000011100011100001111001010100;
        10'd571: TDATA = 37'b0000111001011001000100101111001001101;
        10'd572: TDATA = 37'b0000111010010101101001101111001000110;
        10'd573: TDATA = 37'b0000111011010010001011001111001000000;
        10'd574: TDATA = 37'b0000111100001110101001001111000111001;
        10'd575: TDATA = 37'b0000111101001011000100001111000110010;
        10'd576: TDATA = 37'b0000111110000111011011001111000101011;
        10'd577: TDATA = 37'b0000111111000011101111101111000100101;
        10'd578: TDATA = 37'b0001000000000000000000001111000011110;
        10'd579: TDATA = 37'b0001000000111100001101101111000010111;
        10'd580: TDATA = 37'b0001000001111000010111101111000010001;
        10'd581: TDATA = 37'b0001000010110100011110001111000001010;
        10'd582: TDATA = 37'b0001000011110000100001101111000000100;
        10'd583: TDATA = 37'b0001000100101100100010001110111111101;
        10'd584: TDATA = 37'b0001000101101000011110101110111110110;
        10'd585: TDATA = 37'b0001000110100100011000001110111110000;
        10'd586: TDATA = 37'b0001000111100000001110101110111101001;
        10'd587: TDATA = 37'b0001001000011100000001101110111100011;
        10'd588: TDATA = 37'b0001001001010111110001101110111011100;
        10'd589: TDATA = 37'b0001001010010011011110001110111010110;
        10'd590: TDATA = 37'b0001001011001111000111001110111001111;
        10'd591: TDATA = 37'b0001001100001010101101001110111001001;
        10'd592: TDATA = 37'b0001001101000110010000001110111000010;
        10'd593: TDATA = 37'b0001001110000001101111101110110111100;
        10'd594: TDATA = 37'b0001001110111101001100001110110110110;
        10'd595: TDATA = 37'b0001001111111000100101001110110101111;
        10'd596: TDATA = 37'b0001010000110011111011001110110101001;
        10'd597: TDATA = 37'b0001010001101111001110001110110100010;
        10'd598: TDATA = 37'b0001010010101010011101101110110011100;
        10'd599: TDATA = 37'b0001010011100101101010001110110010110;
        10'd600: TDATA = 37'b0001010100100000110011101110110001111;
        10'd601: TDATA = 37'b0001010101011011111001101110110001001;
        10'd602: TDATA = 37'b0001010110010110111100101110110000011;
        10'd603: TDATA = 37'b0001010111010001111100101110101111101;
        10'd604: TDATA = 37'b0001011000001100111001001110101110110;
        10'd605: TDATA = 37'b0001011001000111110010101110101110000;
        10'd606: TDATA = 37'b0001011010000010101001001110101101010;
        10'd607: TDATA = 37'b0001011010111101011100101110101100100;
        10'd608: TDATA = 37'b0001011011111000001101001110101011101;
        10'd609: TDATA = 37'b0001011100110010111010001110101010111;
        10'd610: TDATA = 37'b0001011101101101100100001110101010001;
        10'd611: TDATA = 37'b0001011110101000001011001110101001011;
        10'd612: TDATA = 37'b0001011111100010101111001110101000101;
        10'd613: TDATA = 37'b0001100000011101010000001110100111111;
        10'd614: TDATA = 37'b0001100001010111101110001110100111001;
        10'd615: TDATA = 37'b0001100010010010001001001110100110011;
        10'd616: TDATA = 37'b0001100011001100100000101110100101101;
        10'd617: TDATA = 37'b0001100100000110110101101110100100110;
        10'd618: TDATA = 37'b0001100101000001000111001110100100000;
        10'd619: TDATA = 37'b0001100101111011010101101110100011010;
        10'd620: TDATA = 37'b0001100110110101100001101110100010100;
        10'd621: TDATA = 37'b0001100111101111101010001110100001110;
        10'd622: TDATA = 37'b0001101000101001110000001110100001000;
        10'd623: TDATA = 37'b0001101001100011110010101110100000010;
        10'd624: TDATA = 37'b0001101010011101110010001110011111100;
        10'd625: TDATA = 37'b0001101011010111101111001110011110111;
        10'd626: TDATA = 37'b0001101100010001101001001110011110001;
        10'd627: TDATA = 37'b0001101101001011011111101110011101011;
        10'd628: TDATA = 37'b0001101110000101010011101110011100101;
        10'd629: TDATA = 37'b0001101110111111000100101110011011111;
        10'd630: TDATA = 37'b0001101111111000110010101110011011001;
        10'd631: TDATA = 37'b0001110000110010011101101110011010011;
        10'd632: TDATA = 37'b0001110001101100000101101110011001101;
        10'd633: TDATA = 37'b0001110010100101101011001110011001000;
        10'd634: TDATA = 37'b0001110011011111001101001110011000010;
        10'd635: TDATA = 37'b0001110100011000101100101110010111100;
        10'd636: TDATA = 37'b0001110101010010001001001110010110110;
        10'd637: TDATA = 37'b0001110110001011100011001110010110000;
        10'd638: TDATA = 37'b0001110111000100111001101110010101011;
        10'd639: TDATA = 37'b0001110111111110001101101110010100101;
        10'd640: TDATA = 37'b0001111000110111011110101110010011111;
        10'd641: TDATA = 37'b0001111001110000101100101110010011001;
        10'd642: TDATA = 37'b0001111010101001111000001110010010100;
        10'd643: TDATA = 37'b0001111011100011000000101110010001110;
        10'd644: TDATA = 37'b0001111100011100000110001110010001000;
        10'd645: TDATA = 37'b0001111101010101001000101110010000011;
        10'd646: TDATA = 37'b0001111110001110001000101110001111101;
        10'd647: TDATA = 37'b0001111111000111000101101110001110111;
        10'd648: TDATA = 37'b0010000000000000000000001110001110010;
        10'd649: TDATA = 37'b0010000000111000110111101110001101100;
        10'd650: TDATA = 37'b0010000001110001101100001110001100111;
        10'd651: TDATA = 37'b0010000010101010011110001110001100001;
        10'd652: TDATA = 37'b0010000011100011001101001110001011011;
        10'd653: TDATA = 37'b0010000100011011111001101110001010110;
        10'd654: TDATA = 37'b0010000101010100100011001110001010000;
        10'd655: TDATA = 37'b0010000110001101001010001110001001011;
        10'd656: TDATA = 37'b0010000111000101101110001110001000101;
        10'd657: TDATA = 37'b0010000111111110001111001110001000000;
        10'd658: TDATA = 37'b0010001000110110101101101110000111010;
        10'd659: TDATA = 37'b0010001001101111001001001110000110101;
        10'd660: TDATA = 37'b0010001010100111100010001110000101111;
        10'd661: TDATA = 37'b0010001011011111111000101110000101010;
        10'd662: TDATA = 37'b0010001100011000001100001110000100100;
        10'd663: TDATA = 37'b0010001101010000011101001110000011111;
        10'd664: TDATA = 37'b0010001110001000101011001110000011010;
        10'd665: TDATA = 37'b0010001111000000110110101110000010100;
        10'd666: TDATA = 37'b0010001111111000111111001110000001111;
        10'd667: TDATA = 37'b0010010000110001000101001110000001001;
        10'd668: TDATA = 37'b0010010001101001001000101110000000100;
        10'd669: TDATA = 37'b0010010010100001001001001101111111111;
        10'd670: TDATA = 37'b0010010011011001000111001101111111001;
        10'd671: TDATA = 37'b0010010100010001000010101101111110100;
        10'd672: TDATA = 37'b0010010101001000111011001101111101111;
        10'd673: TDATA = 37'b0010010110000000110001001101111101001;
        10'd674: TDATA = 37'b0010010110111000100100001101111100100;
        10'd675: TDATA = 37'b0010010111110000010101001101111011111;
        10'd676: TDATA = 37'b0010011000101000000011001101111011001;
        10'd677: TDATA = 37'b0010011001011111101110001101111010100;
        10'd678: TDATA = 37'b0010011010010111010111001101111001111;
        10'd679: TDATA = 37'b0010011011001110111101001101111001010;
        10'd680: TDATA = 37'b0010011100000110100000101101111000100;
        10'd681: TDATA = 37'b0010011100111110000001101101110111111;
        10'd682: TDATA = 37'b0010011101110101011111101101110111010;
        10'd683: TDATA = 37'b0010011110101100111011101101110110101;
        10'd684: TDATA = 37'b0010011111100100010100101101110110000;
        10'd685: TDATA = 37'b0010100000011011101011001101110101010;
        10'd686: TDATA = 37'b0010100001010010111111001101110100101;
        10'd687: TDATA = 37'b0010100010001010010000001101110100000;
        10'd688: TDATA = 37'b0010100011000001011111001101110011011;
        10'd689: TDATA = 37'b0010100011111000101011001101110010110;
        10'd690: TDATA = 37'b0010100100101111110100101101110010001;
        10'd691: TDATA = 37'b0010100101100110111100001101110001100;
        10'd692: TDATA = 37'b0010100110011110000000101101110000110;
        10'd693: TDATA = 37'b0010100111010101000010001101110000001;
        10'd694: TDATA = 37'b0010101000001100000001101101101111100;
        10'd695: TDATA = 37'b0010101001000010111110101101101110111;
        10'd696: TDATA = 37'b0010101001111001111001001101101110010;
        10'd697: TDATA = 37'b0010101010110000110000101101101101101;
        10'd698: TDATA = 37'b0010101011100111100110001101101101000;
        10'd699: TDATA = 37'b0010101100011110011001001101101100011;
        10'd700: TDATA = 37'b0010101101010101001001001101101011110;
        10'd701: TDATA = 37'b0010101110001011110111001101101011001;
        10'd702: TDATA = 37'b0010101111000010100010101101101010100;
        10'd703: TDATA = 37'b0010101111111001001011001101101001111;
        10'd704: TDATA = 37'b0010110000101111110001101101101001010;
        10'd705: TDATA = 37'b0010110001100110010101001101101000101;
        10'd706: TDATA = 37'b0010110010011100110110101101101000000;
        10'd707: TDATA = 37'b0010110011010011010101101101100111011;
        10'd708: TDATA = 37'b0010110100001001110010001101100110110;
        10'd709: TDATA = 37'b0010110101000000001100001101100110001;
        10'd710: TDATA = 37'b0010110101110110100011101101100101101;
        10'd711: TDATA = 37'b0010110110101100111000101101100101000;
        10'd712: TDATA = 37'b0010110111100011001011001101100100011;
        10'd713: TDATA = 37'b0010111000011001011011101101100011110;
        10'd714: TDATA = 37'b0010111001001111101001001101100011001;
        10'd715: TDATA = 37'b0010111010000101110100101101100010100;
        10'd716: TDATA = 37'b0010111010111011111101001101100001111;
        10'd717: TDATA = 37'b0010111011110010000011101101100001011;
        10'd718: TDATA = 37'b0010111100101000001000001101100000110;
        10'd719: TDATA = 37'b0010111101011110001001101101100000001;
        10'd720: TDATA = 37'b0010111110010100001000101101011111100;
        10'd721: TDATA = 37'b0010111111001010000101101101011110111;
        10'd722: TDATA = 37'b0011000000000000000000001101011110011;
        10'd723: TDATA = 37'b0011000000110101111000001101011101110;
        10'd724: TDATA = 37'b0011000001101011101110001101011101001;
        10'd725: TDATA = 37'b0011000010100001100001001101011100100;
        10'd726: TDATA = 37'b0011000011010111010010001101011011111;
        10'd727: TDATA = 37'b0011000100001101000000101101011011011;
        10'd728: TDATA = 37'b0011000101000010101101001101011010110;
        10'd729: TDATA = 37'b0011000101111000010110101101011010001;
        10'd730: TDATA = 37'b0011000110101101111110001101011001101;
        10'd731: TDATA = 37'b0011000111100011100011001101011001000;
        10'd732: TDATA = 37'b0011001000011001000110001101011000011;
        10'd733: TDATA = 37'b0011001001001110100110101101010111111;
        10'd734: TDATA = 37'b0011001010000100000100101101010111010;
        10'd735: TDATA = 37'b0011001010111001100000101101010110101;
        10'd736: TDATA = 37'b0011001011101110111010001101010110001;
        10'd737: TDATA = 37'b0011001100100100010001001101010101100;
        10'd738: TDATA = 37'b0011001101011001100110001101010100111;
        10'd739: TDATA = 37'b0011001110001110111000101101010100011;
        10'd740: TDATA = 37'b0011001111000100001000101101010011110;
        10'd741: TDATA = 37'b0011001111111001010110101101010011010;
        10'd742: TDATA = 37'b0011010000101110100010001101010010101;
        10'd743: TDATA = 37'b0011010001100011101011101101010010000;
        10'd744: TDATA = 37'b0011010010011000110010101101010001100;
        10'd745: TDATA = 37'b0011010011001101110111001101010000111;
        10'd746: TDATA = 37'b0011010100000010111001101101010000011;
        10'd747: TDATA = 37'b0011010100110111111010001101001111110;
        10'd748: TDATA = 37'b0011010101101100110111101101001111010;
        10'd749: TDATA = 37'b0011010110100001110011101101001110101;
        10'd750: TDATA = 37'b0011010111010110101100101101001110001;
        10'd751: TDATA = 37'b0011011000001011100100001101001101100;
        10'd752: TDATA = 37'b0011011001000000011001001101001101000;
        10'd753: TDATA = 37'b0011011001110101001011101101001100011;
        10'd754: TDATA = 37'b0011011010101001111100001101001011111;
        10'd755: TDATA = 37'b0011011011011110101010001101001011010;
        10'd756: TDATA = 37'b0011011100010011010110001101001010110;
        10'd757: TDATA = 37'b0011011101000111111111101101001010001;
        10'd758: TDATA = 37'b0011011101111100100111001101001001101;
        10'd759: TDATA = 37'b0011011110110001001100101101001001000;
        10'd760: TDATA = 37'b0011011111100101101111101101001000100;
        10'd761: TDATA = 37'b0011100000011010010000001101000111111;
        10'd762: TDATA = 37'b0011100001001110101110101101000111011;
        10'd763: TDATA = 37'b0011100010000011001011001101000110111;
        10'd764: TDATA = 37'b0011100010110111100101101101000110010;
        10'd765: TDATA = 37'b0011100011101011111101101101000101110;
        10'd766: TDATA = 37'b0011100100100000010011001101000101001;
        10'd767: TDATA = 37'b0011100101010100100111001101000100101;
        10'd768: TDATA = 37'b0011100110001000111000101101000100001;
        10'd769: TDATA = 37'b0011100110111101000111101101000011100;
        10'd770: TDATA = 37'b0011100111110001010100101101000011000;
        10'd771: TDATA = 37'b0011101000100101011111101101000010100;
        10'd772: TDATA = 37'b0011101001011001101000101101000001111;
        10'd773: TDATA = 37'b0011101010001101101111001101000001011;
        10'd774: TDATA = 37'b0011101011000001110011101101000000111;
        10'd775: TDATA = 37'b0011101011110101110110001101000000010;
        10'd776: TDATA = 37'b0011101100101001110110001100111111110;
        10'd777: TDATA = 37'b0011101101011101110100001100111111010;
        10'd778: TDATA = 37'b0011101110010001110000001100111110110;
        10'd779: TDATA = 37'b0011101111000101101001101100111110001;
        10'd780: TDATA = 37'b0011101111111001100001001100111101101;
        10'd781: TDATA = 37'b0011110000101101010110101100111101001;
        10'd782: TDATA = 37'b0011110001100001001010001100111100101;
        10'd783: TDATA = 37'b0011110010010100111011101100111100000;
        10'd784: TDATA = 37'b0011110011001000101010101100111011100;
        10'd785: TDATA = 37'b0011110011111100010111101100111011000;
        10'd786: TDATA = 37'b0011110100110000000010101100111010100;
        10'd787: TDATA = 37'b0011110101100011101011001100111010000;
        10'd788: TDATA = 37'b0011110110010111010010001100111001011;
        10'd789: TDATA = 37'b0011110111001010110110101100111000111;
        10'd790: TDATA = 37'b0011110111111110011001001100111000011;
        10'd791: TDATA = 37'b0011111000110001111001101100110111111;
        10'd792: TDATA = 37'b0011111001100101010111101100110111011;
        10'd793: TDATA = 37'b0011111010011000110100001100110110110;
        10'd794: TDATA = 37'b0011111011001100001110001100110110010;
        10'd795: TDATA = 37'b0011111011111111100110101100110101110;
        10'd796: TDATA = 37'b0011111100110010111100101100110101010;
        10'd797: TDATA = 37'b0011111101100110010000101100110100110;
        10'd798: TDATA = 37'b0011111110011001100010101100110100010;
        10'd799: TDATA = 37'b0011111111001100110010001100110011110;
        10'd800: TDATA = 37'b0100000000000000000000001100110011010;
        10'd801: TDATA = 37'b0100000000110011001100001100110010110;
        10'd802: TDATA = 37'b0100000001100110010101101100110010001;
        10'd803: TDATA = 37'b0100000010011001011101001100110001101;
        10'd804: TDATA = 37'b0100000011001100100011001100110001001;
        10'd805: TDATA = 37'b0100000011111111100110101100110000101;
        10'd806: TDATA = 37'b0100000100110010101000001100110000001;
        10'd807: TDATA = 37'b0100000101100101100111101100101111101;
        10'd808: TDATA = 37'b0100000110011000100101001100101111001;
        10'd809: TDATA = 37'b0100000111001011100000101100101110101;
        10'd810: TDATA = 37'b0100000111111110011010001100101110001;
        10'd811: TDATA = 37'b0100001000110001010001101100101101101;
        10'd812: TDATA = 37'b0100001001100100000111001100101101001;
        10'd813: TDATA = 37'b0100001010010110111010101100101100101;
        10'd814: TDATA = 37'b0100001011001001101100001100101100001;
        10'd815: TDATA = 37'b0100001011111100011011101100101011101;
        10'd816: TDATA = 37'b0100001100101111001001001100101011001;
        10'd817: TDATA = 37'b0100001101100001110101001100101010101;
        10'd818: TDATA = 37'b0100001110010100011110101100101010001;
        10'd819: TDATA = 37'b0100001111000111000110001100101001101;
        10'd820: TDATA = 37'b0100001111111001101011101100101001001;
        10'd821: TDATA = 37'b0100010000101100001111001100101000101;
        10'd822: TDATA = 37'b0100010001011110110000101100101000001;
        10'd823: TDATA = 37'b0100010010010001010000101100100111101;
        10'd824: TDATA = 37'b0100010011000011101110001100100111001;
        10'd825: TDATA = 37'b0100010011110110001010001100100110110;
        10'd826: TDATA = 37'b0100010100101000100011101100100110010;
        10'd827: TDATA = 37'b0100010101011010111011101100100101110;
        10'd828: TDATA = 37'b0100010110001101010001101100100101010;
        10'd829: TDATA = 37'b0100010110111111100101101100100100110;
        10'd830: TDATA = 37'b0100010111110001110111101100100100010;
        10'd831: TDATA = 37'b0100011000100100000111101100100011110;
        10'd832: TDATA = 37'b0100011001010110010101101100100011010;
        10'd833: TDATA = 37'b0100011010001000100001101100100010110;
        10'd834: TDATA = 37'b0100011010111010101100001100100010011;
        10'd835: TDATA = 37'b0100011011101100110100101100100001111;
        10'd836: TDATA = 37'b0100011100011110111010101100100001011;
        10'd837: TDATA = 37'b0100011101010000111111101100100000111;
        10'd838: TDATA = 37'b0100011110000011000010001100100000011;
        10'd839: TDATA = 37'b0100011110110101000010101100011111111;
        10'd840: TDATA = 37'b0100011111100111000001101100011111100;
        10'd841: TDATA = 37'b0100100000011000111110001100011111000;
        10'd842: TDATA = 37'b0100100001001010111001001100011110100;
        10'd843: TDATA = 37'b0100100001111100110010101100011110000;
        10'd844: TDATA = 37'b0100100010101110101001101100011101100;
        10'd845: TDATA = 37'b0100100011100000011110101100011101001;
        10'd846: TDATA = 37'b0100100100010010010010001100011100101;
        10'd847: TDATA = 37'b0100100101000100000011101100011100001;
        10'd848: TDATA = 37'b0100100101110101110011101100011011101;
        10'd849: TDATA = 37'b0100100110100111100001001100011011010;
        10'd850: TDATA = 37'b0100100111011001001101001100011010110;
        10'd851: TDATA = 37'b0100101000001010110111001100011010010;
        10'd852: TDATA = 37'b0100101000111100011111001100011001110;
        10'd853: TDATA = 37'b0100101001101110000101101100011001011;
        10'd854: TDATA = 37'b0100101010011111101010001100011000111;
        10'd855: TDATA = 37'b0100101011010001001100101100011000011;
        10'd856: TDATA = 37'b0100101100000010101101001100011000000;
        10'd857: TDATA = 37'b0100101100110100001100001100010111100;
        10'd858: TDATA = 37'b0100101101100101101001001100010111000;
        10'd859: TDATA = 37'b0100101110010111000100101100010110101;
        10'd860: TDATA = 37'b0100101111001000011101101100010110001;
        10'd861: TDATA = 37'b0100101111111001110101001100010101101;
        10'd862: TDATA = 37'b0100110000101011001011001100010101010;
        10'd863: TDATA = 37'b0100110001011100011110101100010100110;
        10'd864: TDATA = 37'b0100110010001101110000101100010100010;
        10'd865: TDATA = 37'b0100110010111111000001001100010011111;
        10'd866: TDATA = 37'b0100110011110000001111101100010011011;
        10'd867: TDATA = 37'b0100110100100001011100001100010010111;
        10'd868: TDATA = 37'b0100110101010010100110101100010010100;
        10'd869: TDATA = 37'b0100110110000011101111101100010010000;
        10'd870: TDATA = 37'b0100110110110100110110101100010001100;
        10'd871: TDATA = 37'b0100110111100101111100001100010001001;
        10'd872: TDATA = 37'b0100111000010110111111101100010000101;
        10'd873: TDATA = 37'b0100111001001000000001001100010000010;
        10'd874: TDATA = 37'b0100111001111001000001001100001111110;
        10'd875: TDATA = 37'b0100111010101001111111001100001111010;
        10'd876: TDATA = 37'b0100111011011010111011101100001110111;
        10'd877: TDATA = 37'b0100111100001011110110001100001110011;
        10'd878: TDATA = 37'b0100111100111100101111001100001110000;
        10'd879: TDATA = 37'b0100111101101101100101101100001101100;
        10'd880: TDATA = 37'b0100111110011110011011001100001101001;
        10'd881: TDATA = 37'b0100111111001111001110101100001100101;
        10'd882: TDATA = 37'b0101000000000000000000001100001100010;
        10'd883: TDATA = 37'b0101000000110000110000001100001011110;
        10'd884: TDATA = 37'b0101000001100001011110001100001011010;
        10'd885: TDATA = 37'b0101000010010010001010101100001010111;
        10'd886: TDATA = 37'b0101000011000010110101001100001010011;
        10'd887: TDATA = 37'b0101000011110011011110001100001010000;
        10'd888: TDATA = 37'b0101000100100100000101001100001001100;
        10'd889: TDATA = 37'b0101000101010100101010001100001001001;
        10'd890: TDATA = 37'b0101000110000101001101101100001000101;
        10'd891: TDATA = 37'b0101000110110101101111101100001000010;
        10'd892: TDATA = 37'b0101000111100110001111101100000111110;
        10'd893: TDATA = 37'b0101001000010110101110001100000111011;
        10'd894: TDATA = 37'b0101001001000111001010101100000110111;
        10'd895: TDATA = 37'b0101001001110111100101101100000110100;
        10'd896: TDATA = 37'b0101001010100111111110101100000110001;
        10'd897: TDATA = 37'b0101001011011000010110001100000101101;
        10'd898: TDATA = 37'b0101001100001000101100001100000101010;
        10'd899: TDATA = 37'b0101001100111000111111101100000100110;
        10'd900: TDATA = 37'b0101001101101001010010001100000100011;
        10'd901: TDATA = 37'b0101001110011001100010101100000011111;
        10'd902: TDATA = 37'b0101001111001001110001101100000011100;
        10'd903: TDATA = 37'b0101001111111001111110101100000011001;
        10'd904: TDATA = 37'b0101010000101010001010001100000010101;
        10'd905: TDATA = 37'b0101010001011010010011101100000010010;
        10'd906: TDATA = 37'b0101010010001010011011101100000001110;
        10'd907: TDATA = 37'b0101010010111010100010001100000001011;
        10'd908: TDATA = 37'b0101010011101010100110101100000001000;
        10'd909: TDATA = 37'b0101010100011010101001101100000000100;
        10'd910: TDATA = 37'b0101010101001010101010101100000000001;
        10'd911: TDATA = 37'b0101010101111010101010001011111111101;
        10'd912: TDATA = 37'b0101010110101010101000001011111111010;
        10'd913: TDATA = 37'b0101010111011010100100001011111110111;
        10'd914: TDATA = 37'b0101011000001010011110101011111110011;
        10'd915: TDATA = 37'b0101011000111010010111101011111110000;
        10'd916: TDATA = 37'b0101011001101010001110101011111101101;
        10'd917: TDATA = 37'b0101011010011010000100001011111101001;
        10'd918: TDATA = 37'b0101011011001001111000001011111100110;
        10'd919: TDATA = 37'b0101011011111001101010001011111100011;
        10'd920: TDATA = 37'b0101011100101001011010101011111011111;
        10'd921: TDATA = 37'b0101011101011001001001001011111011100;
        10'd922: TDATA = 37'b0101011110001000110110101011111011001;
        10'd923: TDATA = 37'b0101011110111000100010001011111010101;
        10'd924: TDATA = 37'b0101011111101000001011101011111010010;
        10'd925: TDATA = 37'b0101100000010111110100001011111001111;
        10'd926: TDATA = 37'b0101100001000111011010101011111001011;
        10'd927: TDATA = 37'b0101100001110110111111101011111001000;
        10'd928: TDATA = 37'b0101100010100110100010101011111000101;
        10'd929: TDATA = 37'b0101100011010110000100001011111000010;
        10'd930: TDATA = 37'b0101100100000101100100001011110111110;
        10'd931: TDATA = 37'b0101100100110101000010101011110111011;
        10'd932: TDATA = 37'b0101100101100100011111001011110111000;
        10'd933: TDATA = 37'b0101100110010011111010101011110110101;
        10'd934: TDATA = 37'b0101100111000011010100001011110110001;
        10'd935: TDATA = 37'b0101100111110010101011101011110101110;
        10'd936: TDATA = 37'b0101101000100010000010001011110101011;
        10'd937: TDATA = 37'b0101101001010001010110101011110101000;
        10'd938: TDATA = 37'b0101101010000000101001101011110100100;
        10'd939: TDATA = 37'b0101101010101111111010101011110100001;
        10'd940: TDATA = 37'b0101101011011111001010101011110011110;
        10'd941: TDATA = 37'b0101101100001110011000101011110011011;
        10'd942: TDATA = 37'b0101101100111101100101001011110010111;
        10'd943: TDATA = 37'b0101101101101100110000001011110010100;
        10'd944: TDATA = 37'b0101101110011011111001101011110010001;
        10'd945: TDATA = 37'b0101101111001011000001001011110001110;
        10'd946: TDATA = 37'b0101101111111010000111101011110001011;
        10'd947: TDATA = 37'b0101110000101001001100001011110001000;
        10'd948: TDATA = 37'b0101110001011000001111001011110000100;
        10'd949: TDATA = 37'b0101110010000111010000001011110000001;
        10'd950: TDATA = 37'b0101110010110110010000001011101111110;
        10'd951: TDATA = 37'b0101110011100101001110001011101111011;
        10'd952: TDATA = 37'b0101110100010100001011001011101111000;
        10'd953: TDATA = 37'b0101110101000011000110001011101110101;
        10'd954: TDATA = 37'b0101110101110001111111101011101110001;
        10'd955: TDATA = 37'b0101110110100000110111101011101101110;
        10'd956: TDATA = 37'b0101110111001111101101101011101101011;
        10'd957: TDATA = 37'b0101110111111110100010101011101101000;
        10'd958: TDATA = 37'b0101111000101101010101101011101100101;
        10'd959: TDATA = 37'b0101111001011100000111001011101100010;
        10'd960: TDATA = 37'b0101111010001010110111101011101011111;
        10'd961: TDATA = 37'b0101111010111001100110001011101011011;
        10'd962: TDATA = 37'b0101111011101000010011001011101011000;
        10'd963: TDATA = 37'b0101111100010110111110001011101010101;
        10'd964: TDATA = 37'b0101111101000101101000001011101010010;
        10'd965: TDATA = 37'b0101111101110100010000101011101001111;
        10'd966: TDATA = 37'b0101111110100010110111001011101001100;
        10'd967: TDATA = 37'b0101111111010001011100101011101001001;
        10'd968: TDATA = 37'b0110000000000000000000001011101000110;
        10'd969: TDATA = 37'b0110000000101110100010001011101000011;
        10'd970: TDATA = 37'b0110000001011101000010101011101000000;
        10'd971: TDATA = 37'b0110000010001011100010001011100111101;
        10'd972: TDATA = 37'b0110000010111001111111101011100111010;
        10'd973: TDATA = 37'b0110000011101000011011101011100110110;
        10'd974: TDATA = 37'b0110000100010110110110001011100110011;
        10'd975: TDATA = 37'b0110000101000101001111001011100110000;
        10'd976: TDATA = 37'b0110000101110011100110001011100101101;
        10'd977: TDATA = 37'b0110000110100001111100001011100101010;
        10'd978: TDATA = 37'b0110000111010000010000101011100100111;
        10'd979: TDATA = 37'b0110000111111110100011101011100100100;
        10'd980: TDATA = 37'b0110001000101100110101001011100100001;
        10'd981: TDATA = 37'b0110001001011011000100101011100011110;
        10'd982: TDATA = 37'b0110001010001001010011001011100011011;
        10'd983: TDATA = 37'b0110001010110111100000001011100011000;
        10'd984: TDATA = 37'b0110001011100101101011001011100010101;
        10'd985: TDATA = 37'b0110001100010011110101001011100010010;
        10'd986: TDATA = 37'b0110001101000001111101101011100001111;
        10'd987: TDATA = 37'b0110001101110000000100001011100001100;
        10'd988: TDATA = 37'b0110001110011110001001101011100001001;
        10'd989: TDATA = 37'b0110001111001100001101101011100000110;
        10'd990: TDATA = 37'b0110001111111010010000001011100000011;
        10'd991: TDATA = 37'b0110010000101000010000101011100000000;
        10'd992: TDATA = 37'b0110010001010110010000001011011111101;
        10'd993: TDATA = 37'b0110010010000100001110001011011111010;
        10'd994: TDATA = 37'b0110010010110010001010101011011110111;
        10'd995: TDATA = 37'b0110010011100000000101101011011110100;
        10'd996: TDATA = 37'b0110010100001101111111001011011110001;
        10'd997: TDATA = 37'b0110010100111011110111001011011101111;
        10'd998: TDATA = 37'b0110010101101001101101101011011101100;
        10'd999: TDATA = 37'b0110010110010111100010101011011101001;
        10'd1000: TDATA = 37'b0110010111000101010110001011011100110;
        10'd1001: TDATA = 37'b0110010111110011001000001011011100011;
        10'd1002: TDATA = 37'b0110011000100000111001001011011100000;
        10'd1003: TDATA = 37'b0110011001001110101000001011011011101;
        10'd1004: TDATA = 37'b0110011001111100010110001011011011010;
        10'd1005: TDATA = 37'b0110011010101010000010001011011010111;
        10'd1006: TDATA = 37'b0110011011010111101101001011011010100;
        10'd1007: TDATA = 37'b0110011100000101010110101011011010001;
        10'd1008: TDATA = 37'b0110011100110010111110001011011001110;
        10'd1009: TDATA = 37'b0110011101100000100100101011011001100;
        10'd1010: TDATA = 37'b0110011110001110001001101011011001001;
        10'd1011: TDATA = 37'b0110011110111011101101101011011000110;
        10'd1012: TDATA = 37'b0110011111101001001111101011011000011;
        10'd1013: TDATA = 37'b0110100000010110110000001011011000000;
        10'd1014: TDATA = 37'b0110100001000100001111101011010111101;
        10'd1015: TDATA = 37'b0110100001110001101101101011010111010;
        10'd1016: TDATA = 37'b0110100010011111001001101011010110111;
        10'd1017: TDATA = 37'b0110100011001100100100101011010110101;
        10'd1018: TDATA = 37'b0110100011111001111110001011010110010;
        10'd1019: TDATA = 37'b0110100100100111010110101011010101111;
        10'd1020: TDATA = 37'b0110100101010100101101001011010101100;
        10'd1021: TDATA = 37'b0110100110000010000010101011010101001;
        10'd1022: TDATA = 37'b0110100110101111010110001011010100110;
        10'd1023: TDATA = 37'b0110100111011100101000101011010100011;
        10'd0: TDATA = 37'b0110101000001001111001110110101000001;
        10'd1: TDATA = 37'b0110101001100100010111110110100110110;
        10'd2: TDATA = 37'b0110101010111110101111110110100101011;
        10'd3: TDATA = 37'b0110101100011001000010010110100011111;
        10'd4: TDATA = 37'b0110101101110011001111010110100010100;
        10'd5: TDATA = 37'b0110101111001101010110110110100001001;
        10'd6: TDATA = 37'b0110110000100111011000010110011111110;
        10'd7: TDATA = 37'b0110110010000001010100110110011110011;
        10'd8: TDATA = 37'b0110110011011011001011010110011101000;
        10'd9: TDATA = 37'b0110110100110100111100010110011011101;
        10'd10: TDATA = 37'b0110110110001110100111110110011010010;
        10'd11: TDATA = 37'b0110110111101000001110010110011000111;
        10'd12: TDATA = 37'b0110111001000001101110110110010111100;
        10'd13: TDATA = 37'b0110111010011011001001110110010110001;
        10'd14: TDATA = 37'b0110111011110100011111110110010100110;
        10'd15: TDATA = 37'b0110111101001101101111110110010011011;
        10'd16: TDATA = 37'b0110111110100110111010110110010010000;
        10'd17: TDATA = 37'b0111000000000000000000010110010000110;
        10'd18: TDATA = 37'b0111000001011001000000010110001111011;
        10'd19: TDATA = 37'b0111000010110001111011010110001110000;
        10'd20: TDATA = 37'b0111000100001010110000010110001100101;
        10'd21: TDATA = 37'b0111000101100011100000010110001011011;
        10'd22: TDATA = 37'b0111000110111100001011010110001010000;
        10'd23: TDATA = 37'b0111001000010100110000110110001000101;
        10'd24: TDATA = 37'b0111001001101101010000110110000111011;
        10'd25: TDATA = 37'b0111001011000101101011010110000110000;
        10'd26: TDATA = 37'b0111001100011110000000110110000100110;
        10'd27: TDATA = 37'b0111001101110110010001010110000011011;
        10'd28: TDATA = 37'b0111001111001110011100010110000010001;
        10'd29: TDATA = 37'b0111010000100110100010010110000000110;
        10'd30: TDATA = 37'b0111010001111110100010110101111111100;
        10'd31: TDATA = 37'b0111010011010110011110010101111110010;
        10'd32: TDATA = 37'b0111010100101110010100010101111100111;
        10'd33: TDATA = 37'b0111010110000110000101110101111011101;
        10'd34: TDATA = 37'b0111010111011101110001010101111010011;
        10'd35: TDATA = 37'b0111011000110101011000010101111001000;
        10'd36: TDATA = 37'b0111011010001100111001110101110111110;
        10'd37: TDATA = 37'b0111011011100100010110110101110110100;
        10'd38: TDATA = 37'b0111011100111011101101110101110101010;
        10'd39: TDATA = 37'b0111011110010011000000010101110100000;
        10'd40: TDATA = 37'b0111011111101010001101110101110010110;
        10'd41: TDATA = 37'b0111100001000001010101110101110001011;
        10'd42: TDATA = 37'b0111100010011000011001010101110000001;
        10'd43: TDATA = 37'b0111100011101111010111010101101110111;
        10'd44: TDATA = 37'b0111100101000110010000110101101101101;
        10'd45: TDATA = 37'b0111100110011101000100110101101100011;
        10'd46: TDATA = 37'b0111100111110011110100010101101011001;
        10'd47: TDATA = 37'b0111101001001010011110010101101010000;
        10'd48: TDATA = 37'b0111101010100001000011110101101000110;
        10'd49: TDATA = 37'b0111101011110111100011110101100111100;
        10'd50: TDATA = 37'b0111101101001101111111010101100110010;
        10'd51: TDATA = 37'b0111101110100100010101110101100101000;
        10'd52: TDATA = 37'b0111101111111010100111010101100011110;
        10'd53: TDATA = 37'b0111110001010000110011110101100010100;
        10'd54: TDATA = 37'b0111110010100110111011110101100001011;
        10'd55: TDATA = 37'b0111110011111100111110110101100000001;
        10'd56: TDATA = 37'b0111110101010010111100110101011110111;
        10'd57: TDATA = 37'b0111110110101000110110010101011101110;
        10'd58: TDATA = 37'b0111110111111110101010010101011100100;
        10'd59: TDATA = 37'b0111111001010100011010010101011011010;
        10'd60: TDATA = 37'b0111111010101010000100110101011010001;
        10'd61: TDATA = 37'b0111111011111111101010110101011000111;
        10'd62: TDATA = 37'b0111111101010101001100010101010111110;
        10'd63: TDATA = 37'b0111111110101010101000110101010110100;
        10'd64: TDATA = 37'b1000000000000000000000010101010101011;
        10'd65: TDATA = 37'b1000000001010101010011010101010100001;
        10'd66: TDATA = 37'b1000000010101010100001010101010011000;
        10'd67: TDATA = 37'b1000000011111111101010110101010001110;
        10'd68: TDATA = 37'b1000000101010100101111110101010000101;
        10'd69: TDATA = 37'b1000000110101001101111110101001111100;
        10'd70: TDATA = 37'b1000000111111110101011010101001110010;
        10'd71: TDATA = 37'b1000001001010011100010010101001101001;
        10'd72: TDATA = 37'b1000001010101000010100010101001100000;
        10'd73: TDATA = 37'b1000001011111101000001110101001010110;
        10'd74: TDATA = 37'b1000001101010001101010110101001001101;
        10'd75: TDATA = 37'b1000001110100110001110110101001000100;
        10'd76: TDATA = 37'b1000001111111010101110010101000111011;
        10'd77: TDATA = 37'b1000010001001111001001010101000110001;
        10'd78: TDATA = 37'b1000010010100011011111110101000101000;
        10'd79: TDATA = 37'b1000010011110111110001110101000011111;
        10'd80: TDATA = 37'b1000010101001011111111010101000010110;
        10'd81: TDATA = 37'b1000010110100000000111110101000001101;
        10'd82: TDATA = 37'b1000010111110100001100010101000000100;
        10'd83: TDATA = 37'b1000011001001000001011110100111111011;
        10'd84: TDATA = 37'b1000011010011100000110110100111110010;
        10'd85: TDATA = 37'b1000011011101111111101110100111101001;
        10'd86: TDATA = 37'b1000011101000011101111110100111100000;
        10'd87: TDATA = 37'b1000011110010111011101010100111010111;
        10'd88: TDATA = 37'b1000011111101011000110110100111001110;
        10'd89: TDATA = 37'b1000100000111110101011010100111000101;
        10'd90: TDATA = 37'b1000100010010010001011110100110111100;
        10'd91: TDATA = 37'b1000100011100101100111110100110110011;
        10'd92: TDATA = 37'b1000100100111000111111010100110101010;
        10'd93: TDATA = 37'b1000100110001100010010010100110100010;
        10'd94: TDATA = 37'b1000100111011111100000110100110011001;
        10'd95: TDATA = 37'b1000101000110010101010110100110010000;
        10'd96: TDATA = 37'b1000101010000101110000110100110000111;
        10'd97: TDATA = 37'b1000101011011000110010010100101111111;
        10'd98: TDATA = 37'b1000101100101011101111010100101110110;
        10'd99: TDATA = 37'b1000101101111110101000010100101101101;
        10'd100: TDATA = 37'b1000101111010001011100110100101100101;
        10'd101: TDATA = 37'b1000110000100100001100110100101011100;
        10'd102: TDATA = 37'b1000110001110110111000110100101010011;
        10'd103: TDATA = 37'b1000110011001001100000010100101001011;
        10'd104: TDATA = 37'b1000110100011100000011010100101000010;
        10'd105: TDATA = 37'b1000110101101110100010010100100111010;
        10'd106: TDATA = 37'b1000110111000000111100110100100110001;
        10'd107: TDATA = 37'b1000111000010011010011010100100101000;
        10'd108: TDATA = 37'b1000111001100101100101010100100100000;
        10'd109: TDATA = 37'b1000111010110111110011010100100010111;
        10'd110: TDATA = 37'b1000111100001001111100110100100001111;
        10'd111: TDATA = 37'b1000111101011100000010010100100000111;
        10'd112: TDATA = 37'b1000111110101110000011010100011111110;
        10'd113: TDATA = 37'b1001000000000000000000010100011110110;
        10'd114: TDATA = 37'b1001000001010001111001010100011101101;
        10'd115: TDATA = 37'b1001000010100011101101110100011100101;
        10'd116: TDATA = 37'b1001000011110101011110010100011011101;
        10'd117: TDATA = 37'b1001000101000111001010010100011010100;
        10'd118: TDATA = 37'b1001000110011000110010010100011001100;
        10'd119: TDATA = 37'b1001000111101010010110010100011000100;
        10'd120: TDATA = 37'b1001001000111011110110010100010111100;
        10'd121: TDATA = 37'b1001001010001101010001110100010110011;
        10'd122: TDATA = 37'b1001001011011110101001110100010101011;
        10'd123: TDATA = 37'b1001001100101111111100110100010100011;
        10'd124: TDATA = 37'b1001001110000001001100010100010011011;
        10'd125: TDATA = 37'b1001001111010010010111110100010010011;
        10'd126: TDATA = 37'b1001010000100011011110110100010001010;
        10'd127: TDATA = 37'b1001010001110100100010010100010000010;
        10'd128: TDATA = 37'b1001010011000101100001010100001111010;
        10'd129: TDATA = 37'b1001010100010110011100010100001110010;
        10'd130: TDATA = 37'b1001010101100111010011010100001101010;
        10'd131: TDATA = 37'b1001010110111000000110010100001100010;
        10'd132: TDATA = 37'b1001011000001000110101010100001011010;
        10'd133: TDATA = 37'b1001011001011001100000010100001010010;
        10'd134: TDATA = 37'b1001011010101010000111010100001001010;
        10'd135: TDATA = 37'b1001011011111010101010010100001000010;
        10'd136: TDATA = 37'b1001011101001011001001010100000111010;
        10'd137: TDATA = 37'b1001011110011011100100010100000110010;
        10'd138: TDATA = 37'b1001011111101011111011010100000101010;
        10'd139: TDATA = 37'b1001100000111100001110010100000100010;
        10'd140: TDATA = 37'b1001100010001100011101010100000011010;
        10'd141: TDATA = 37'b1001100011011100101000110100000010010;
        10'd142: TDATA = 37'b1001100100101100101111110100000001011;
        10'd143: TDATA = 37'b1001100101111100110011010100000000011;
        10'd144: TDATA = 37'b1001100111001100110010110011111111011;
        10'd145: TDATA = 37'b1001101000011100101110010011111110011;
        10'd146: TDATA = 37'b1001101001101100100101110011111101011;
        10'd147: TDATA = 37'b1001101010111100011001110011111100100;
        10'd148: TDATA = 37'b1001101100001100001001110011111011100;
        10'd149: TDATA = 37'b1001101101011011110101110011111010100;
        10'd150: TDATA = 37'b1001101110101011011101110011111001101;
        10'd151: TDATA = 37'b1001101111111011000010010011111000101;
        10'd152: TDATA = 37'b1001110001001010100010110011110111101;
        10'd153: TDATA = 37'b1001110010011001111111010011110110110;
        10'd154: TDATA = 37'b1001110011101001011000010011110101110;
        10'd155: TDATA = 37'b1001110100111000101101010011110100110;
        10'd156: TDATA = 37'b1001110110000111111110010011110011111;
        10'd157: TDATA = 37'b1001110111010111001011110011110010111;
        10'd158: TDATA = 37'b1001111000100110010101010011110010000;
        10'd159: TDATA = 37'b1001111001110101011011010011110001000;
        10'd160: TDATA = 37'b1001111011000100011101010011110000000;
        10'd161: TDATA = 37'b1001111100010011011011110011101111001;
        10'd162: TDATA = 37'b1001111101100010010110010011101110001;
        10'd163: TDATA = 37'b1001111110110001001101010011101101010;
        10'd164: TDATA = 37'b1010000000000000000000010011101100010;
        10'd165: TDATA = 37'b1010000001001110101111110011101011011;
        10'd166: TDATA = 37'b1010000010011101011011010011101010100;
        10'd167: TDATA = 37'b1010000011101100000011010011101001100;
        10'd168: TDATA = 37'b1010000100111010100111010011101000101;
        10'd169: TDATA = 37'b1010000110001001000111110011100111101;
        10'd170: TDATA = 37'b1010000111010111100100110011100110110;
        10'd171: TDATA = 37'b1010001000100101111101110011100101111;
        10'd172: TDATA = 37'b1010001001110100010011010011100100111;
        10'd173: TDATA = 37'b1010001011000010100101010011100100000;
        10'd174: TDATA = 37'b1010001100010000110011010011100011001;
        10'd175: TDATA = 37'b1010001101011110111110010011100010001;
        10'd176: TDATA = 37'b1010001110101101000100110011100001010;
        10'd177: TDATA = 37'b1010001111111011001000010011100000011;
        10'd178: TDATA = 37'b1010010001001001000111110011011111100;
        10'd179: TDATA = 37'b1010010010010111000011110011011110100;
        10'd180: TDATA = 37'b1010010011100100111100010011011101101;
        10'd181: TDATA = 37'b1010010100110010110001010011011100110;
        10'd182: TDATA = 37'b1010010110000000100010010011011011111;
        10'd183: TDATA = 37'b1010010111001110001111110011011011000;
        10'd184: TDATA = 37'b1010011000011011111001110011011010001;
        10'd185: TDATA = 37'b1010011001101001100000010011011001001;
        10'd186: TDATA = 37'b1010011010110111000011010011011000010;
        10'd187: TDATA = 37'b1010011100000100100010110011010111011;
        10'd188: TDATA = 37'b1010011101010001111110110011010110100;
        10'd189: TDATA = 37'b1010011110011111010110110011010101101;
        10'd190: TDATA = 37'b1010011111101100101011110011010100110;
        10'd191: TDATA = 37'b1010100000111001111100110011010011111;
        10'd192: TDATA = 37'b1010100010000111001010110011010011000;
        10'd193: TDATA = 37'b1010100011010100010100110011010010001;
        10'd194: TDATA = 37'b1010100100100001011011010011010001010;
        10'd195: TDATA = 37'b1010100101101110011110110011010000011;
        10'd196: TDATA = 37'b1010100110111011011110010011001111100;
        10'd197: TDATA = 37'b1010101000001000011010110011001110101;
        10'd198: TDATA = 37'b1010101001010101010011010011001101110;
        10'd199: TDATA = 37'b1010101010100010001000110011001100111;
        10'd200: TDATA = 37'b1010101011101110111010110011001100000;
        10'd201: TDATA = 37'b1010101100111011101001010011001011001;
        10'd202: TDATA = 37'b1010101110001000010011110011001010010;
        10'd203: TDATA = 37'b1010101111010100111011110011001001100;
        10'd204: TDATA = 37'b1010110000100001011111110011001000101;
        10'd205: TDATA = 37'b1010110001101110000000010011000111110;
        10'd206: TDATA = 37'b1010110010111010011101110011000110111;
        10'd207: TDATA = 37'b1010110100000110110111010011000110000;
        10'd208: TDATA = 37'b1010110101010011001101110011000101010;
        10'd209: TDATA = 37'b1010110110011111100000110011000100011;
        10'd210: TDATA = 37'b1010110111101011110000110011000011100;
        10'd211: TDATA = 37'b1010111000110111111100110011000010101;
        10'd212: TDATA = 37'b1010111010000100000101110011000001111;
        10'd213: TDATA = 37'b1010111011010000001011010011000001000;
        10'd214: TDATA = 37'b1010111100011100001101110011000000001;
        10'd215: TDATA = 37'b1010111101101000001100110010111111010;
        10'd216: TDATA = 37'b1010111110110100001000010010111110100;
        10'd217: TDATA = 37'b1011000000000000000000010010111101101;
        10'd218: TDATA = 37'b1011000001001011110101010010111100110;
        10'd219: TDATA = 37'b1011000010010111100110110010111100000;
        10'd220: TDATA = 37'b1011000011100011010100110010111011001;
        10'd221: TDATA = 37'b1011000100101110111111110010111010011;
        10'd222: TDATA = 37'b1011000101111010100111010010111001100;
        10'd223: TDATA = 37'b1011000111000110001011110010111000101;
        10'd224: TDATA = 37'b1011001000010001101100110010110111111;
        10'd225: TDATA = 37'b1011001001011101001010010010110111000;
        10'd226: TDATA = 37'b1011001010101000100100110010110110010;
        10'd227: TDATA = 37'b1011001011110011111100010010110101011;
        10'd228: TDATA = 37'b1011001100111111010000010010110100101;
        10'd229: TDATA = 37'b1011001110001010100000110010110011110;
        10'd230: TDATA = 37'b1011001111010101101110010010110011000;
        10'd231: TDATA = 37'b1011010000100000111000010010110010001;
        10'd232: TDATA = 37'b1011010001101011111111010010110001011;
        10'd233: TDATA = 37'b1011010010110111000010110010110000100;
        10'd234: TDATA = 37'b1011010100000010000011010010101111110;
        10'd235: TDATA = 37'b1011010101001101000000110010101110111;
        10'd236: TDATA = 37'b1011010110010111111010110010101110001;
        10'd237: TDATA = 37'b1011010111100010110001110010101101011;
        10'd238: TDATA = 37'b1011011000101101100101010010101100100;
        10'd239: TDATA = 37'b1011011001111000010101110010101011110;
        10'd240: TDATA = 37'b1011011011000011000011010010101010111;
        10'd241: TDATA = 37'b1011011100001101101101010010101010001;
        10'd242: TDATA = 37'b1011011101011000010100010010101001011;
        10'd243: TDATA = 37'b1011011110100010110111110010101000100;
        10'd244: TDATA = 37'b1011011111101101011000110010100111110;
        10'd245: TDATA = 37'b1011100000110111110110010010100111000;
        10'd246: TDATA = 37'b1011100010000010010000010010100110001;
        10'd247: TDATA = 37'b1011100011001100100111110010100101011;
        10'd248: TDATA = 37'b1011100100010110111011110010100100101;
        10'd249: TDATA = 37'b1011100101100001001100110010100011111;
        10'd250: TDATA = 37'b1011100110101011011010010010100011000;
        10'd251: TDATA = 37'b1011100111110101100100110010100010010;
        10'd252: TDATA = 37'b1011101000111111101100110010100001100;
        10'd253: TDATA = 37'b1011101010001001110001010010100000110;
        10'd254: TDATA = 37'b1011101011010011110010010010100000000;
        10'd255: TDATA = 37'b1011101100011101110000110010011111001;
        10'd256: TDATA = 37'b1011101101100111101011110010011110011;
        10'd257: TDATA = 37'b1011101110110001100011110010011101101;
        10'd258: TDATA = 37'b1011101111111011011001010010011100111;
        10'd259: TDATA = 37'b1011110001000101001011010010011100001;
        10'd260: TDATA = 37'b1011110010001110111001110010011011011;
        10'd261: TDATA = 37'b1011110011011000100101110010011010101;
        10'd262: TDATA = 37'b1011110100100010001110110010011001111;
        10'd263: TDATA = 37'b1011110101101011110100010010011001000;
        10'd264: TDATA = 37'b1011110110110101010111010010011000010;
        10'd265: TDATA = 37'b1011110111111110110110110010010111100;
        10'd266: TDATA = 37'b1011111001001000010011010010010110110;
        10'd267: TDATA = 37'b1011111010010001101101010010010110000;
        10'd268: TDATA = 37'b1011111011011011000011110010010101010;
        10'd269: TDATA = 37'b1011111100100100010111010010010100100;
        10'd270: TDATA = 37'b1011111101101101100111110010010011110;
        10'd271: TDATA = 37'b1011111110110110110101110010010011000;
        10'd272: TDATA = 37'b1100000000000000000000010010010010010;
        10'd273: TDATA = 37'b1100000001001001000111110010010001100;
        10'd274: TDATA = 37'b1100000010010010001100110010010000110;
        10'd275: TDATA = 37'b1100000011011011001110010010010000000;
        10'd276: TDATA = 37'b1100000100100100001100110010001111010;
        10'd277: TDATA = 37'b1100000101101101001000110010001110101;
        10'd278: TDATA = 37'b1100000110110110000001110010001101111;
        10'd279: TDATA = 37'b1100000111111110110111010010001101001;
        10'd280: TDATA = 37'b1100001001000111101010010010001100011;
        10'd281: TDATA = 37'b1100001010010000011010010010001011101;
        10'd282: TDATA = 37'b1100001011011001000111010010001010111;
        10'd283: TDATA = 37'b1100001100100001110001010010001010001;
        10'd284: TDATA = 37'b1100001101101010011000110010001001011;
        10'd285: TDATA = 37'b1100001110110010111100110010001000110;
        10'd286: TDATA = 37'b1100001111111011011110010010001000000;
        10'd287: TDATA = 37'b1100010001000011111100110010000111010;
        10'd288: TDATA = 37'b1100010010001100011000010010000110100;
        10'd289: TDATA = 37'b1100010011010100110000110010000101110;
        10'd290: TDATA = 37'b1100010100011101000110110010000101001;
        10'd291: TDATA = 37'b1100010101100101011001110010000100011;
        10'd292: TDATA = 37'b1100010110101101101001110010000011101;
        10'd293: TDATA = 37'b1100010111110101110110110010000010111;
        10'd294: TDATA = 37'b1100011000111110000000110010000010010;
        10'd295: TDATA = 37'b1100011010000110001000010010000001100;
        10'd296: TDATA = 37'b1100011011001110001100110010000000110;
        10'd297: TDATA = 37'b1100011100010110001110010010000000000;
        10'd298: TDATA = 37'b1100011101011110001101010001111111011;
        10'd299: TDATA = 37'b1100011110100110001001010001111110101;
        10'd300: TDATA = 37'b1100011111101110000010010001111101111;
        10'd301: TDATA = 37'b1100100000110101111000110001111101010;
        10'd302: TDATA = 37'b1100100001111101101100010001111100100;
        10'd303: TDATA = 37'b1100100011000101011100110001111011111;
        10'd304: TDATA = 37'b1100100100001101001010110001111011001;
        10'd305: TDATA = 37'b1100100101010100110101110001111010011;
        10'd306: TDATA = 37'b1100100110011100011101110001111001110;
        10'd307: TDATA = 37'b1100100111100100000011010001111001000;
        10'd308: TDATA = 37'b1100101000101011100110010001111000010;
        10'd309: TDATA = 37'b1100101001110011000101110001110111101;
        10'd310: TDATA = 37'b1100101010111010100010110001110110111;
        10'd311: TDATA = 37'b1100101100000001111101010001110110010;
        10'd312: TDATA = 37'b1100101101001001010100110001110101100;
        10'd313: TDATA = 37'b1100101110010000101001010001110100111;
        10'd314: TDATA = 37'b1100101111010111111011010001110100001;
        10'd315: TDATA = 37'b1100110000011111001010110001110011100;
        10'd316: TDATA = 37'b1100110001100110010111010001110010110;
        10'd317: TDATA = 37'b1100110010101101100000110001110010001;
        10'd318: TDATA = 37'b1100110011110100100111110001110001011;
        10'd319: TDATA = 37'b1100110100111011101011110001110000110;
        10'd320: TDATA = 37'b1100110110000010101101010001110000000;
        10'd321: TDATA = 37'b1100110111001001101100010001101111011;
        10'd322: TDATA = 37'b1100111000010000101000010001101110101;
        10'd323: TDATA = 37'b1100111001010111100001010001101110000;
        10'd324: TDATA = 37'b1100111010011110010111110001101101010;
        10'd325: TDATA = 37'b1100111011100101001011110001101100101;
        10'd326: TDATA = 37'b1100111100101011111100110001101100000;
        10'd327: TDATA = 37'b1100111101110010101011010001101011010;
        10'd328: TDATA = 37'b1100111110111001010111010001101010101;
        10'd329: TDATA = 37'b1101000000000000000000010001101001111;
        10'd330: TDATA = 37'b1101000001000110100110110001101001010;
        10'd331: TDATA = 37'b1101000010001101001010010001101000101;
        10'd332: TDATA = 37'b1101000011010011101011010001100111111;
        10'd333: TDATA = 37'b1101000100011010001001110001100111010;
        10'd334: TDATA = 37'b1101000101100000100101010001100110101;
        10'd335: TDATA = 37'b1101000110100110111110010001100101111;
        10'd336: TDATA = 37'b1101000111101101010100110001100101010;
        10'd337: TDATA = 37'b1101001000110011101000010001100100101;
        10'd338: TDATA = 37'b1101001001111001111001110001100011111;
        10'd339: TDATA = 37'b1101001011000000000111110001100011010;
        10'd340: TDATA = 37'b1101001100000110010011110001100010101;
        10'd341: TDATA = 37'b1101001101001100011100110001100010000;
        10'd342: TDATA = 37'b1101001110010010100011010001100001010;
        10'd343: TDATA = 37'b1101001111011000100111010001100000101;
        10'd344: TDATA = 37'b1101010000011110101000010001100000000;
        10'd345: TDATA = 37'b1101010001100100100111010001011111011;
        10'd346: TDATA = 37'b1101010010101010100011010001011110101;
        10'd347: TDATA = 37'b1101010011110000011100110001011110000;
        10'd348: TDATA = 37'b1101010100110110010011010001011101011;
        10'd349: TDATA = 37'b1101010101111100000111110001011100110;
        10'd350: TDATA = 37'b1101010111000001111001010001011100001;
        10'd351: TDATA = 37'b1101011000000111101000010001011011011;
        10'd352: TDATA = 37'b1101011001001101010100110001011010110;
        10'd353: TDATA = 37'b1101011010010010111110110001011010001;
        10'd354: TDATA = 37'b1101011011011000100101110001011001100;
        10'd355: TDATA = 37'b1101011100011110001010110001011000111;
        10'd356: TDATA = 37'b1101011101100011101100110001011000010;
        10'd357: TDATA = 37'b1101011110101001001100010001010111101;
        10'd358: TDATA = 37'b1101011111101110101001010001010111000;
        10'd359: TDATA = 37'b1101100000110100000011110001010110010;
        10'd360: TDATA = 37'b1101100001111001011011110001010101101;
        10'd361: TDATA = 37'b1101100010111110110001010001010101000;
        10'd362: TDATA = 37'b1101100100000100000100010001010100011;
        10'd363: TDATA = 37'b1101100101001001010100010001010011110;
        10'd364: TDATA = 37'b1101100110001110100010010001010011001;
        10'd365: TDATA = 37'b1101100111010011101101010001010010100;
        10'd366: TDATA = 37'b1101101000011000110110010001010001111;
        10'd367: TDATA = 37'b1101101001011101111100010001010001010;
        10'd368: TDATA = 37'b1101101010100010111111110001010000101;
        10'd369: TDATA = 37'b1101101011101000000001010001010000000;
        10'd370: TDATA = 37'b1101101100101100111111110001001111011;
        10'd371: TDATA = 37'b1101101101110001111100010001001110110;
        10'd372: TDATA = 37'b1101101110110110110101110001001110001;
        10'd373: TDATA = 37'b1101101111111011101100110001001101100;
        10'd374: TDATA = 37'b1101110001000000100001110001001100111;
        10'd375: TDATA = 37'b1101110010000101010011110001001100010;
        10'd376: TDATA = 37'b1101110011001010000011110001001011101;
        10'd377: TDATA = 37'b1101110100001110110000110001001011000;
        10'd378: TDATA = 37'b1101110101010011011011110001001010011;
        10'd379: TDATA = 37'b1101110110011000000011110001001001110;
        10'd380: TDATA = 37'b1101110111011100101001110001001001001;
        10'd381: TDATA = 37'b1101111000100001001101010001001000100;
        10'd382: TDATA = 37'b1101111001100101101110010001000111111;
        10'd383: TDATA = 37'b1101111010101010001100010001000111011;
        10'd384: TDATA = 37'b1101111011101110101000110001000110110;
        10'd385: TDATA = 37'b1101111100110011000010010001000110001;
        10'd386: TDATA = 37'b1101111101110111011001010001000101100;
        10'd387: TDATA = 37'b1101111110111011101101110001000100111;
        10'd388: TDATA = 37'b1110000000000000000000010001000100010;
        10'd389: TDATA = 37'b1110000001000100010000010001000011101;
        10'd390: TDATA = 37'b1110000010001000011101110001000011000;
        10'd391: TDATA = 37'b1110000011001100101000110001000010100;
        10'd392: TDATA = 37'b1110000100010000110001010001000001111;
        10'd393: TDATA = 37'b1110000101010100110111010001000001010;
        10'd394: TDATA = 37'b1110000110011000111011010001000000101;
        10'd395: TDATA = 37'b1110000111011100111100010001000000000;
        10'd396: TDATA = 37'b1110001000100000111011010000111111100;
        10'd397: TDATA = 37'b1110001001100100111000010000111110111;
        10'd398: TDATA = 37'b1110001010101000110010010000111110010;
        10'd399: TDATA = 37'b1110001011101100101010010000111101101;
        10'd400: TDATA = 37'b1110001100110000011111010000111101000;
        10'd401: TDATA = 37'b1110001101110100010010010000111100100;
        10'd402: TDATA = 37'b1110001110111000000011010000111011111;
        10'd403: TDATA = 37'b1110001111111011110001010000111011010;
        10'd404: TDATA = 37'b1110010000111111011101010000111010101;
        10'd405: TDATA = 37'b1110010010000011000110110000111010001;
        10'd406: TDATA = 37'b1110010011000110101110010000111001100;
        10'd407: TDATA = 37'b1110010100001010010010110000111000111;
        10'd408: TDATA = 37'b1110010101001101110101010000111000011;
        10'd409: TDATA = 37'b1110010110010001010101110000110111110;
        10'd410: TDATA = 37'b1110010111010100110011010000110111001;
        10'd411: TDATA = 37'b1110011000011000001110110000110110101;
        10'd412: TDATA = 37'b1110011001011011100111110000110110000;
        10'd413: TDATA = 37'b1110011010011110111110110000110101011;
        10'd414: TDATA = 37'b1110011011100010010011010000110100111;
        10'd415: TDATA = 37'b1110011100100101100101010000110100010;
        10'd416: TDATA = 37'b1110011101101000110101010000110011101;
        10'd417: TDATA = 37'b1110011110101100000010110000110011001;
        10'd418: TDATA = 37'b1110011111101111001101110000110010100;
        10'd419: TDATA = 37'b1110100000110010010110110000110001111;
        10'd420: TDATA = 37'b1110100001110101011101010000110001011;
        10'd421: TDATA = 37'b1110100010111000100001010000110000110;
        10'd422: TDATA = 37'b1110100011111011100011010000110000010;
        10'd423: TDATA = 37'b1110100100111110100011010000101111101;
        10'd424: TDATA = 37'b1110100110000001100000010000101111000;
        10'd425: TDATA = 37'b1110100111000100011011110000101110100;
        10'd426: TDATA = 37'b1110101000000111010100010000101101111;
        10'd427: TDATA = 37'b1110101001001010001010110000101101011;
        10'd428: TDATA = 37'b1110101010001100111111010000101100110;
        10'd429: TDATA = 37'b1110101011001111110001010000101100010;
        10'd430: TDATA = 37'b1110101100010010100000110000101011101;
        10'd431: TDATA = 37'b1110101101010101001110010000101011001;
        10'd432: TDATA = 37'b1110101110010111111001010000101010100;
        10'd433: TDATA = 37'b1110101111011010100010010000101010000;
        10'd434: TDATA = 37'b1110110000011101001000110000101001011;
        10'd435: TDATA = 37'b1110110001011111101101010000101000111;
        10'd436: TDATA = 37'b1110110010100010001111010000101000010;
        10'd437: TDATA = 37'b1110110011100100101111010000100111110;
        10'd438: TDATA = 37'b1110110100100111001100110000100111001;
        10'd439: TDATA = 37'b1110110101101001101000010000100110101;
        10'd440: TDATA = 37'b1110110110101100000001110000100110000;
        10'd441: TDATA = 37'b1110110111101110011000110000100101100;
        10'd442: TDATA = 37'b1110111000110000101101010000100100111;
        10'd443: TDATA = 37'b1110111001110010111111110000100100011;
        10'd444: TDATA = 37'b1110111010110101010000010000100011110;
        10'd445: TDATA = 37'b1110111011110111011110010000100011010;
        10'd446: TDATA = 37'b1110111100111001101001110000100010101;
        10'd447: TDATA = 37'b1110111101111011110011110000100010001;
        10'd448: TDATA = 37'b1110111110111101111011010000100001101;
        10'd449: TDATA = 37'b1111000000000000000000010000100001000;
        10'd450: TDATA = 37'b1111000001000010000011010000100000100;
        10'd451: TDATA = 37'b1111000010000100000100010000011111111;
        10'd452: TDATA = 37'b1111000011000110000010110000011111011;
        10'd453: TDATA = 37'b1111000100000111111111010000011110111;
        10'd454: TDATA = 37'b1111000101001001111001010000011110010;
        10'd455: TDATA = 37'b1111000110001011110001110000011101110;
        10'd456: TDATA = 37'b1111000111001101100111010000011101010;
        10'd457: TDATA = 37'b1111001000001111011011010000011100101;
        10'd458: TDATA = 37'b1111001001010001001100110000011100001;
        10'd459: TDATA = 37'b1111001010010010111100010000011011101;
        10'd460: TDATA = 37'b1111001011010100101001010000011011000;
        10'd461: TDATA = 37'b1111001100010110010100010000011010100;
        10'd462: TDATA = 37'b1111001101010111111101010000011010000;
        10'd463: TDATA = 37'b1111001110011001100100010000011001011;
        10'd464: TDATA = 37'b1111001111011011001000110000011000111;
        10'd465: TDATA = 37'b1111010000011100101011010000011000011;
        10'd466: TDATA = 37'b1111010001011110001011010000010111110;
        10'd467: TDATA = 37'b1111010010011111101001010000010111010;
        10'd468: TDATA = 37'b1111010011100001000101110000010110110;
        10'd469: TDATA = 37'b1111010100100010011111010000010110010;
        10'd470: TDATA = 37'b1111010101100011110111010000010101101;
        10'd471: TDATA = 37'b1111010110100101001100110000010101001;
        10'd472: TDATA = 37'b1111010111100110100000010000010100101;
        10'd473: TDATA = 37'b1111011000100111110001110000010100001;
        10'd474: TDATA = 37'b1111011001101001000000110000010011100;
        10'd475: TDATA = 37'b1111011010101010001101110000010011000;
        10'd476: TDATA = 37'b1111011011101011011000110000010010100;
        10'd477: TDATA = 37'b1111011100101100100001110000010010000;
        10'd478: TDATA = 37'b1111011101101101101000110000010001011;
        10'd479: TDATA = 37'b1111011110101110101101010000010000111;
        10'd480: TDATA = 37'b1111011111101111101111110000010000011;
        10'd481: TDATA = 37'b1111100000110000110000010000001111111;
        10'd482: TDATA = 37'b1111100001110001101110110000001111011;
        10'd483: TDATA = 37'b1111100010110010101011010000001110111;
        10'd484: TDATA = 37'b1111100011110011100101010000001110010;
        10'd485: TDATA = 37'b1111100100110100011101010000001101110;
        10'd486: TDATA = 37'b1111100101110101010011110000001101010;
        10'd487: TDATA = 37'b1111100110110110000111110000001100110;
        10'd488: TDATA = 37'b1111100111110110111001010000001100010;
        10'd489: TDATA = 37'b1111101000110111101001010000001011110;
        10'd490: TDATA = 37'b1111101001111000010110110000001011001;
        10'd491: TDATA = 37'b1111101010111001000010110000001010101;
        10'd492: TDATA = 37'b1111101011111001101100010000001010001;
        10'd493: TDATA = 37'b1111101100111010010011110000001001101;
        10'd494: TDATA = 37'b1111101101111010111001010000001001001;
        10'd495: TDATA = 37'b1111101110111011011100110000001000101;
        10'd496: TDATA = 37'b1111101111111011111110010000001000001;
        10'd497: TDATA = 37'b1111110000111100011101110000000111101;
        10'd498: TDATA = 37'b1111110001111100111010110000000111001;
        10'd499: TDATA = 37'b1111110010111101010110010000000110101;
        10'd500: TDATA = 37'b1111110011111101101111010000000110000;
        10'd501: TDATA = 37'b1111110100111110000110110000000101100;
        10'd502: TDATA = 37'b1111110101111110011011110000000101000;
        10'd503: TDATA = 37'b1111110110111110101110110000000100100;
        10'd504: TDATA = 37'b1111110111111110111111110000000100000;
        10'd505: TDATA = 37'b1111111000111111001111010000000011100;
        10'd506: TDATA = 37'b1111111001111111011100010000000011000;
        10'd507: TDATA = 37'b1111111010111111100111010000000010100;
        10'd508: TDATA = 37'b1111111011111111110000010000000010000;
        10'd509: TDATA = 37'b1111111100111111110111010000000001100;
        10'd510: TDATA = 37'b1111111101111111111100010000000001000;
        10'd511: TDATA = 37'b1111111110111111111111010000000000100;
        endcase
    end
    endfunction

    wire [7:0] ex;
    assign ex = x[30:23];
    
    wire [9:0] key;
    wire [13:0] h;
    assign key = x[23:14];
    assign h = x[13:0];

    wire [36:0] tdata;
    assign tdata = TDATA(key);

    wire [22:0] rtx0;
    wire [13:0] rtx0_inv;
    assign rtx0 = tdata[36:14];
    assign rtx0_inv = tdata[13:0];

    wire check_zero;
    assign check_zero = (x[30:0] == 31'b0);

    wire [7:0] ey;
    assign ey = (check_zero) ? 8'b0: 8'd63 + ex[7:1] + ex[0] + (x[23:2] == {1'b0,{21{1'b1}}} & x[1:0] != 2'b0);

    wire [36:0] my_extend;
    assign my_extend = {rtx0,14'b0} + rtx0_inv * h;

    wire [22:0] my;
    assign my = (check_zero) ? 23'b0: my_extend[36:14];

    assign y = {1'b0,ey,my};

endmodule

