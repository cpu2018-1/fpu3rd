module finv(
    input wire [31:0] x,
    output wire [31:0] y
);

    function [37:0] TDATA (
	input [10:0] ML
    );
    begin
        casex(ML)
        11'd0: TDATA = 38'b00000000000000000000000100000000000000;
        11'd1: TDATA = 38'b11111111110000000000100011111111110000;
        11'd2: TDATA = 38'b11111111100000000010000011111111100000;
        11'd3: TDATA = 38'b11111111010000000100100011111111010000;
        11'd4: TDATA = 38'b11111111000000001000000011111111000000;
        11'd5: TDATA = 38'b11111110110000001100100011111110110000;
        11'd6: TDATA = 38'b11111110100000010010000011111110100000;
        11'd7: TDATA = 38'b11111110010000011000011011111110010000;
        11'd8: TDATA = 38'b11111110000000011111111011111110000000;
        11'd9: TDATA = 38'b11111101110000101000011011111101110000;
        11'd10: TDATA = 38'b11111101100000110001110011111101100000;
        11'd11: TDATA = 38'b11111101010000111100001011111101010000;
        11'd12: TDATA = 38'b11111101000001000111101011111101000001;
        11'd13: TDATA = 38'b11111100110001010100000011111100110001;
        11'd14: TDATA = 38'b11111100100001100001011011111100100001;
        11'd15: TDATA = 38'b11111100010001101111101011111100010001;
        11'd16: TDATA = 38'b11111100000001111111000011111100000001;
        11'd17: TDATA = 38'b11111011110010001111010011111011110100;
        11'd18: TDATA = 38'b11111011100010100000101011111011100100;
        11'd19: TDATA = 38'b11111011010010110010111011111011010100;
        11'd20: TDATA = 38'b11111011000011000110001011111011000100;
        11'd21: TDATA = 38'b11111010110011011010010011111010110100;
        11'd22: TDATA = 38'b11111010100011101111011011111010100100;
        11'd23: TDATA = 38'b11111010010100000101101011111010010111;
        11'd24: TDATA = 38'b11111010000100011100101011111010000111;
        11'd25: TDATA = 38'b11111001110100110100110011111001110111;
        11'd26: TDATA = 38'b11111001100101001101110011111001101000;
        11'd27: TDATA = 38'b11111001010101100111110011111001011000;
        11'd28: TDATA = 38'b11111001000110000010110011111001001000;
        11'd29: TDATA = 38'b11111000110110011110101011111000111001;
        11'd30: TDATA = 38'b11111000100110111011100011111000101001;
        11'd31: TDATA = 38'b11111000010111011001011011111000011011;
        11'd32: TDATA = 38'b11111000000111111000001011111000001011;
        11'd33: TDATA = 38'b11110111111000010111111011110111111100;
        11'd34: TDATA = 38'b11110111101000111000100011110111101100;
        11'd35: TDATA = 38'b11110111011001011010010011110111011101;
        11'd36: TDATA = 38'b11110111001001111100110011110111001101;
        11'd37: TDATA = 38'b11110110111010100000011011110111000000;
        11'd38: TDATA = 38'b11110110101011000100111011110110110000;
        11'd39: TDATA = 38'b11110110011011101010010011110110100000;
        11'd40: TDATA = 38'b11110110001100010000101011110110010011;
        11'd41: TDATA = 38'b11110101111100111000000011110110000011;
        11'd42: TDATA = 38'b11110101101101100000010011110101110100;
        11'd43: TDATA = 38'b11110101011110001001100011110101100100;
        11'd44: TDATA = 38'b11110101001110110011101011110101010101;
        11'd45: TDATA = 38'b11110100111111011110110011110101000111;
        11'd46: TDATA = 38'b11110100110000001010110011110100111000;
        11'd47: TDATA = 38'b11110100100000110111110011110100101000;
        11'd48: TDATA = 38'b11110100010001100101101011110100011001;
        11'd49: TDATA = 38'b11110100000010010100100011110100001011;
        11'd50: TDATA = 38'b11110011110011000100010011110011111100;
        11'd51: TDATA = 38'b11110011100011110100111011110011101100;
        11'd52: TDATA = 38'b11110011010100100110100011110011011111;
        11'd53: TDATA = 38'b11110011000101011001001011110011010000;
        11'd54: TDATA = 38'b11110010110110001100100011110011000000;
        11'd55: TDATA = 38'b11110010100111000001000011110010110011;
        11'd56: TDATA = 38'b11110010010111110110010011110010100011;
        11'd57: TDATA = 38'b11110010001000101100100011110010010100;
        11'd58: TDATA = 38'b11110001111001100011101011110010000101;
        11'd59: TDATA = 38'b11110001101010011011110011110001110111;
        11'd60: TDATA = 38'b11110001011011010100110011110001101000;
        11'd61: TDATA = 38'b11110001001100001110110011110001011001;
        11'd62: TDATA = 38'b11110000111101001001100011110001001100;
        11'd63: TDATA = 38'b11110000101110000101010011110000111100;
        11'd64: TDATA = 38'b11110000011111000010000011110000101111;
        11'd65: TDATA = 38'b11110000001111111111100011110000011111;
        11'd66: TDATA = 38'b11110000000000111110000011110000010000;
        11'd67: TDATA = 38'b11101111110001111101011011110000000001;
        11'd68: TDATA = 38'b11101111100010111101110011101111110011;
        11'd69: TDATA = 38'b11101111010011111110111011101111100100;
        11'd70: TDATA = 38'b11101111000101000001000011101111010111;
        11'd71: TDATA = 38'b11101110110110000100000011101111001000;
        11'd72: TDATA = 38'b11101110100111001000000011101110111001;
        11'd73: TDATA = 38'b11101110011000001100110011101110101100;
        11'd74: TDATA = 38'b11101110001001010010100011101110011100;
        11'd75: TDATA = 38'b11101101111010011001001011101110001111;
        11'd76: TDATA = 38'b11101101101011100000101011101110000000;
        11'd77: TDATA = 38'b11101101011100101001001011101101110001;
        11'd78: TDATA = 38'b11101101001101110010011011101101100100;
        11'd79: TDATA = 38'b11101100111110111100101011101101010100;
        11'd80: TDATA = 38'b11101100110000000111110011101101001000;
        11'd81: TDATA = 38'b11101100100001010011110011101100111000;
        11'd82: TDATA = 38'b11101100010010100000101011101100101011;
        11'd83: TDATA = 38'b11101100000011101110011011101100011100;
        11'd84: TDATA = 38'b11101011110100111101000011101100001101;
        11'd85: TDATA = 38'b11101011100110001100100011101100000000;
        11'd86: TDATA = 38'b11101011010111011101000011101011110001;
        11'd87: TDATA = 38'b11101011001000101110010011101011100100;
        11'd88: TDATA = 38'b11101010111010000000100011101011010101;
        11'd89: TDATA = 38'b11101010101011010011100011101011001000;
        11'd90: TDATA = 38'b11101010011100100111100011101010111001;
        11'd91: TDATA = 38'b11101010001101111100011011101010101011;
        11'd92: TDATA = 38'b11101001111111010010001011101010011101;
        11'd93: TDATA = 38'b11101001110000101000101011101010001111;
        11'd94: TDATA = 38'b11101001100010000000001011101010000001;
        11'd95: TDATA = 38'b11101001010011011000100011101001110100;
        11'd96: TDATA = 38'b11101001000100110001101011101001100100;
        11'd97: TDATA = 38'b11101000110110001011110011101001011000;
        11'd98: TDATA = 38'b11101000100111100110110011101001001001;
        11'd99: TDATA = 38'b11101000011001000010100011101000111100;
        11'd100: TDATA = 38'b11101000001010011111010011101000101101;
        11'd101: TDATA = 38'b11100111111011111100110011101000100000;
        11'd102: TDATA = 38'b11100111101101011011010011101000010001;
        11'd103: TDATA = 38'b11100111011110111010100011101000000100;
        11'd104: TDATA = 38'b11100111010000011010101011100111110111;
        11'd105: TDATA = 38'b11100111000001111011101011100111101000;
        11'd106: TDATA = 38'b11100110110011011101100011100111011011;
        11'd107: TDATA = 38'b11100110100101000000010011100111001101;
        11'd108: TDATA = 38'b11100110010110100011111011100111000000;
        11'd109: TDATA = 38'b11100110001000001000010011100110110001;
        11'd110: TDATA = 38'b11100101111001101101101011100110100100;
        11'd111: TDATA = 38'b11100101101011010011110011100110010111;
        11'd112: TDATA = 38'b11100101011100111010110011100110001000;
        11'd113: TDATA = 38'b11100101001110100010101011100101111011;
        11'd114: TDATA = 38'b11100101000000001011011011100101101101;
        11'd115: TDATA = 38'b11100100110001110100111011100101100000;
        11'd116: TDATA = 38'b11100100100011011111011011100101010011;
        11'd117: TDATA = 38'b11100100010101001010101011100101000100;
        11'd118: TDATA = 38'b11100100000110110110110011100100110111;
        11'd119: TDATA = 38'b11100011111000100011101011100100101001;
        11'd120: TDATA = 38'b11100011101010010001100011100100011100;
        11'd121: TDATA = 38'b11100011011100000000001011100100001111;
        11'd122: TDATA = 38'b11100011001101101111101011100100000000;
        11'd123: TDATA = 38'b11100010111111011111111011100011110100;
        11'd124: TDATA = 38'b11100010110001010001001011100011100111;
        11'd125: TDATA = 38'b11100010100011000011001011100011011001;
        11'd126: TDATA = 38'b11100010010100110101111011100011001100;
        11'd127: TDATA = 38'b11100010000110101001101011100010111101;
        11'd128: TDATA = 38'b11100001111000011110001011100010110000;
        11'd129: TDATA = 38'b11100001101010010011100011100010100100;
        11'd130: TDATA = 38'b11100001011100001001101011100010010111;
        11'd131: TDATA = 38'b11100001001110000000101011100010001001;
        11'd132: TDATA = 38'b11100000111111111000100011100001111100;
        11'd133: TDATA = 38'b11100000110001110001001011100001101101;
        11'd134: TDATA = 38'b11100000100011101010101011100001100000;
        11'd135: TDATA = 38'b11100000010101100101000011100001010100;
        11'd136: TDATA = 38'b11100000000111100000001011100001000111;
        11'd137: TDATA = 38'b11011111111001011100001011100000111001;
        11'd138: TDATA = 38'b11011111101011011000111011100000101100;
        11'd139: TDATA = 38'b11011111011101010110100011100000100000;
        11'd140: TDATA = 38'b11011111001111010101000011100000010011;
        11'd141: TDATA = 38'b11011111000001010100010011100000000100;
        11'd142: TDATA = 38'b11011110110011010100010011011111111000;
        11'd143: TDATA = 38'b11011110100101010101001011011111101011;
        11'd144: TDATA = 38'b11011110010111010110111011011111011101;
        11'd145: TDATA = 38'b11011110001001011001011011011111010000;
        11'd146: TDATA = 38'b11011101111011011100110011011111000100;
        11'd147: TDATA = 38'b11011101101101100000111011011110110111;
        11'd148: TDATA = 38'b11011101011111100101111011011110101001;
        11'd149: TDATA = 38'b11011101010001101011101011011110011100;
        11'd150: TDATA = 38'b11011101000011110010010011011110010000;
        11'd151: TDATA = 38'b11011100110101111001101011011110000011;
        11'd152: TDATA = 38'b11011100101000000001111011011101110111;
        11'd153: TDATA = 38'b11011100011010001010111011011101101001;
        11'd154: TDATA = 38'b11011100001100010100110011011101011100;
        11'd155: TDATA = 38'b11011011111110011111011011011101010000;
        11'd156: TDATA = 38'b11011011110000101010110011011101000011;
        11'd157: TDATA = 38'b11011011100010110111000011011100110101;
        11'd158: TDATA = 38'b11011011010101000100000011011100101001;
        11'd159: TDATA = 38'b11011011000111010001111011011100011100;
        11'd160: TDATA = 38'b11011010111001100000100011011100010000;
        11'd161: TDATA = 38'b11011010101011101111111011011100000011;
        11'd162: TDATA = 38'b11011010011110000000001011011011110111;
        11'd163: TDATA = 38'b11011010010000010001001011011011101001;
        11'd164: TDATA = 38'b11011010000010100011000011011011011100;
        11'd165: TDATA = 38'b11011001110100110101100011011011010000;
        11'd166: TDATA = 38'b11011001100111001001000011011011000100;
        11'd167: TDATA = 38'b11011001011001011101001011011010110111;
        11'd168: TDATA = 38'b11011001001011110010001011011010101001;
        11'd169: TDATA = 38'b11011000111110000111111011011010011101;
        11'd170: TDATA = 38'b11011000110000011110100011011010010000;
        11'd171: TDATA = 38'b11011000100010110101111011011010000100;
        11'd172: TDATA = 38'b11011000010101001110000011011001111000;
        11'd173: TDATA = 38'b11011000000111100110111011011001101011;
        11'd174: TDATA = 38'b11010111111010000000101011011001011111;
        11'd175: TDATA = 38'b11010111101100011011001011011001010001;
        11'd176: TDATA = 38'b11010111011110110110011011011001000100;
        11'd177: TDATA = 38'b11010111010001010010011011011000111000;
        11'd178: TDATA = 38'b11010111000011101111010011011000101100;
        11'd179: TDATA = 38'b11010110110110001100111011011000100000;
        11'd180: TDATA = 38'b11010110101000101011010011011000010011;
        11'd181: TDATA = 38'b11010110011011001010011011011000001000;
        11'd182: TDATA = 38'b11010110001101101010010011010111111011;
        11'd183: TDATA = 38'b11010110000000001011000011010111101111;
        11'd184: TDATA = 38'b11010101110010101100100011010111100001;
        11'd185: TDATA = 38'b11010101100101001110110011010111010101;
        11'd186: TDATA = 38'b11010101010111110001110011010111001000;
        11'd187: TDATA = 38'b11010101001010010101101011010110111100;
        11'd188: TDATA = 38'b11010100111100111010001011010110110000;
        11'd189: TDATA = 38'b11010100101111011111100011010110100100;
        11'd190: TDATA = 38'b11010100100010000101101011010110011000;
        11'd191: TDATA = 38'b11010100010100101100100011010110001100;
        11'd192: TDATA = 38'b11010100000111010100001011010110000000;
        11'd193: TDATA = 38'b11010011111001111100100011010101110011;
        11'd194: TDATA = 38'b11010011101100100101101011010101100111;
        11'd195: TDATA = 38'b11010011011111001111101011010101011011;
        11'd196: TDATA = 38'b11010011010001111010010011010101001111;
        11'd197: TDATA = 38'b11010011000100100101110011010101000011;
        11'd198: TDATA = 38'b11010010110111010010000011010100110111;
        11'd199: TDATA = 38'b11010010101001111110111011010100101001;
        11'd200: TDATA = 38'b11010010011100101100101011010100011101;
        11'd201: TDATA = 38'b11010010001111011011001011010100010001;
        11'd202: TDATA = 38'b11010010000010001010011011010100000111;
        11'd203: TDATA = 38'b11010001110100111010011011010011111001;
        11'd204: TDATA = 38'b11010001100111101011001011010011101101;
        11'd205: TDATA = 38'b11010001011010011100101011010011100001;
        11'd206: TDATA = 38'b11010001001101001110111011010011010101;
        11'd207: TDATA = 38'b11010001000000000001111011010011001011;
        11'd208: TDATA = 38'b11010000110010110101100011010010111101;
        11'd209: TDATA = 38'b11010000100101101010000011010010110001;
        11'd210: TDATA = 38'b11010000011000011111010011010010100101;
        11'd211: TDATA = 38'b11010000001011010101010011010010011001;
        11'd212: TDATA = 38'b11001111111110001100000011010010001111;
        11'd213: TDATA = 38'b11001111110001000011100011010010000011;
        11'd214: TDATA = 38'b11001111100011111011110011010001110101;
        11'd215: TDATA = 38'b11001111010110110100101011010001101001;
        11'd216: TDATA = 38'b11001111001001101110011011010001011111;
        11'd217: TDATA = 38'b11001110111100101000110011010001010011;
        11'd218: TDATA = 38'b11001110101111100100000011010001000111;
        11'd219: TDATA = 38'b11001110100010011111111011010000111011;
        11'd220: TDATA = 38'b11001110010101011100100011010000110000;
        11'd221: TDATA = 38'b11001110001000011010000011010000100100;
        11'd222: TDATA = 38'b11001101111011011000001011010000011000;
        11'd223: TDATA = 38'b11001101101110010111000011010000001100;
        11'd224: TDATA = 38'b11001101100001010110100011010000000000;
        11'd225: TDATA = 38'b11001101010100010110111011001111110100;
        11'd226: TDATA = 38'b11001101000111010111111011001111101000;
        11'd227: TDATA = 38'b11001100111010011001110011001111011101;
        11'd228: TDATA = 38'b11001100101101011100010011001111010001;
        11'd229: TDATA = 38'b11001100100000011111100011001111000101;
        11'd230: TDATA = 38'b11001100010011100011100011001110111011;
        11'd231: TDATA = 38'b11001100000110101000001011001110101111;
        11'd232: TDATA = 38'b11001011111001101101101011001110100011;
        11'd233: TDATA = 38'b11001011101100110011110011001110011000;
        11'd234: TDATA = 38'b11001011011111111010101011001110001100;
        11'd235: TDATA = 38'b11001011010011000010010011001110000000;
        11'd236: TDATA = 38'b11001011000110001010100011001101110100;
        11'd237: TDATA = 38'b11001010111001010011101011001101101001;
        11'd238: TDATA = 38'b11001010101100011101011011001101011101;
        11'd239: TDATA = 38'b11001010011111100111111011001101010001;
        11'd240: TDATA = 38'b11001010010010110011000011001101000111;
        11'd241: TDATA = 38'b11001010000101111111000011001100111011;
        11'd242: TDATA = 38'b11001001111001001011101011001100110000;
        11'd243: TDATA = 38'b11001001101100011000111011001100100100;
        11'd244: TDATA = 38'b11001001011111100111000011001100011000;
        11'd245: TDATA = 38'b11001001010010110101110011001100001101;
        11'd246: TDATA = 38'b11001001000110000101010011001100000011;
        11'd247: TDATA = 38'b11001000111001010101100011001011110111;
        11'd248: TDATA = 38'b11001000101100100110011011001011101100;
        11'd249: TDATA = 38'b11001000011111111000000011001011100000;
        11'd250: TDATA = 38'b11001000010011001010010011001011010100;
        11'd251: TDATA = 38'b11001000000110011101011011001011001001;
        11'd252: TDATA = 38'b11000111111001110001001011001010111101;
        11'd253: TDATA = 38'b11000111101101000101100011001010110100;
        11'd254: TDATA = 38'b11000111100000011010110011001010101000;
        11'd255: TDATA = 38'b11000111010011110000100011001010011100;
        11'd256: TDATA = 38'b11000111000111000111001011001010010001;
        11'd257: TDATA = 38'b11000110111010011110011011001010000101;
        11'd258: TDATA = 38'b11000110101101110110011011001001111011;
        11'd259: TDATA = 38'b11000110100001001111000011001001110000;
        11'd260: TDATA = 38'b11000110010100101000011011001001100100;
        11'd261: TDATA = 38'b11000110001000000010100011001001011001;
        11'd262: TDATA = 38'b11000101111011011101010011001001001101;
        11'd263: TDATA = 38'b11000101101110111000101011001001000011;
        11'd264: TDATA = 38'b11000101100010010100111011001000111000;
        11'd265: TDATA = 38'b11000101010101110001101011001000101100;
        11'd266: TDATA = 38'b11000101001001001111010011001000100001;
        11'd267: TDATA = 38'b11000100111100101101100011001000010111;
        11'd268: TDATA = 38'b11000100110000001100011011001000001100;
        11'd269: TDATA = 38'b11000100100011101100000011001000000000;
        11'd270: TDATA = 38'b11000100010111001100011011000111110101;
        11'd271: TDATA = 38'b11000100001010101101011011000111101001;
        11'd272: TDATA = 38'b11000011111110001111000011000111100000;
        11'd273: TDATA = 38'b11000011110001110001011011000111010100;
        11'd274: TDATA = 38'b11000011100101010100100011000111001001;
        11'd275: TDATA = 38'b11000011011000111000010011000110111101;
        11'd276: TDATA = 38'b11000011001100011100101011000110110100;
        11'd277: TDATA = 38'b11000011000000000001110011000110101000;
        11'd278: TDATA = 38'b11000010110011100111101011000110011101;
        11'd279: TDATA = 38'b11000010100111001110000011000110010011;
        11'd280: TDATA = 38'b11000010011010110101010011000110001000;
        11'd281: TDATA = 38'b11000010001110011101001011000101111100;
        11'd282: TDATA = 38'b11000010000010000101101011000101110011;
        11'd283: TDATA = 38'b11000001110101101110111011000101100111;
        11'd284: TDATA = 38'b11000001101001011000110011000101011100;
        11'd285: TDATA = 38'b11000001011101000011010011000101010001;
        11'd286: TDATA = 38'b11000001010000101110100011000101000111;
        11'd287: TDATA = 38'b11000001000100011010011011000100111100;
        11'd288: TDATA = 38'b11000000111000000111000011000100110001;
        11'd289: TDATA = 38'b11000000101011110100010011000100100101;
        11'd290: TDATA = 38'b11000000011111100010010011000100011100;
        11'd291: TDATA = 38'b11000000010011010000111011000100010000;
        11'd292: TDATA = 38'b11000000000111000000001011000100000111;
        11'd293: TDATA = 38'b10111111111010110000000011000011111011;
        11'd294: TDATA = 38'b10111111101110100000101011000011110000;
        11'd295: TDATA = 38'b10111111100010010010000011000011100101;
        11'd296: TDATA = 38'b10111111010110000011111011000011011100;
        11'd297: TDATA = 38'b10111111001001110110100011000011010000;
        11'd298: TDATA = 38'b10111110111101101001111011000011000101;
        11'd299: TDATA = 38'b10111110110001011101110011000010111011;
        11'd300: TDATA = 38'b10111110100101010010011011000010110000;
        11'd301: TDATA = 38'b10111110011001000111110011000010100111;
        11'd302: TDATA = 38'b10111110001100111101101011000010011011;
        11'd303: TDATA = 38'b10111110000000110100010011000010010000;
        11'd304: TDATA = 38'b10111101110100101011100011000010000101;
        11'd305: TDATA = 38'b10111101101000100011100011000001111100;
        11'd306: TDATA = 38'b10111101011100011100000011000001110000;
        11'd307: TDATA = 38'b10111101010000010101010011000001100111;
        11'd308: TDATA = 38'b10111101000100001111010011000001011100;
        11'd309: TDATA = 38'b10111100111000001001110011000001010001;
        11'd310: TDATA = 38'b10111100101100000101000011000001001000;
        11'd311: TDATA = 38'b10111100100000000000111011000000111100;
        11'd312: TDATA = 38'b10111100010011111101011011000000110001;
        11'd313: TDATA = 38'b10111100000111111010101011000000101000;
        11'd314: TDATA = 38'b10111011111011111000011011000000011100;
        11'd315: TDATA = 38'b10111011101111110110111011000000010011;
        11'd316: TDATA = 38'b10111011100011110110000011000000001000;
        11'd317: TDATA = 38'b10111011010111110101111010111111111101;
        11'd318: TDATA = 38'b10111011001011110110010010111111110100;
        11'd319: TDATA = 38'b10111010111111110111011010111111101000;
        11'd320: TDATA = 38'b10111010110011111001001010111111011111;
        11'd321: TDATA = 38'b10111010100111111011100010111111010100;
        11'd322: TDATA = 38'b10111010011011111110100010111111001001;
        11'd323: TDATA = 38'b10111010010000000010001010111111000000;
        11'd324: TDATA = 38'b10111010000100000110100010111110110101;
        11'd325: TDATA = 38'b10111001111000001011011010111110101100;
        11'd326: TDATA = 38'b10111001101100010001000010111110100000;
        11'd327: TDATA = 38'b10111001100000010111010010111110010111;
        11'd328: TDATA = 38'b10111001010100011110001010111110001100;
        11'd329: TDATA = 38'b10111001001000100101110010111110000001;
        11'd330: TDATA = 38'b10111000111100101101111010111101111000;
        11'd331: TDATA = 38'b10111000110000110110101010111101101101;
        11'd332: TDATA = 38'b10111000100101000000001010111101100100;
        11'd333: TDATA = 38'b10111000011001001010001010111101011001;
        11'd334: TDATA = 38'b10111000001101010100111010111101010000;
        11'd335: TDATA = 38'b10111000000001100000010010111101000100;
        11'd336: TDATA = 38'b10110111110101101100010010111100111011;
        11'd337: TDATA = 38'b10110111101001111000111010111100110000;
        11'd338: TDATA = 38'b10110111011110000110001010111100100111;
        11'd339: TDATA = 38'b10110111010010010100000010111100011100;
        11'd340: TDATA = 38'b10110111000110100010100010111100010011;
        11'd341: TDATA = 38'b10110110111010110001101010111100001000;
        11'd342: TDATA = 38'b10110110101111000001100010111011111111;
        11'd343: TDATA = 38'b10110110100011010001111010111011110100;
        11'd344: TDATA = 38'b10110110010111100010111010111011101001;
        11'd345: TDATA = 38'b10110110001011110100100010111011100000;
        11'd346: TDATA = 38'b10110110000000000110111010111011010111;
        11'd347: TDATA = 38'b10110101110100011001110010111011001100;
        11'd348: TDATA = 38'b10110101101000101101010010111011000001;
        11'd349: TDATA = 38'b10110101011101000001100010111010111000;
        11'd350: TDATA = 38'b10110101010001010110010010111010101111;
        11'd351: TDATA = 38'b10110101000101101011101010111010100100;
        11'd352: TDATA = 38'b10110100111010000001110010111010011011;
        11'd353: TDATA = 38'b10110100101110011000011010111010010000;
        11'd354: TDATA = 38'b10110100100010101111101010111010000101;
        11'd355: TDATA = 38'b10110100010111000111100010111001111100;
        11'd356: TDATA = 38'b10110100001011100000000010111001110011;
        11'd357: TDATA = 38'b10110011111111111001010010111001101000;
        11'd358: TDATA = 38'b10110011110100010011000010111001011111;
        11'd359: TDATA = 38'b10110011101000101101010010111001010100;
        11'd360: TDATA = 38'b10110011011101001000010010111001001100;
        11'd361: TDATA = 38'b10110011010001100011111010111001000001;
        11'd362: TDATA = 38'b10110011000110000000001010111000111000;
        11'd363: TDATA = 38'b10110010111010011100111010111000101101;
        11'd364: TDATA = 38'b10110010101110111010011010111000100100;
        11'd365: TDATA = 38'b10110010100011011000011010111000011001;
        11'd366: TDATA = 38'b10110010010111110111001010111000010000;
        11'd367: TDATA = 38'b10110010001100010110011010111000000111;
        11'd368: TDATA = 38'b10110010000000110110010010110111111100;
        11'd369: TDATA = 38'b10110001110101010110110010110111110011;
        11'd370: TDATA = 38'b10110001101001110111111010110111101000;
        11'd371: TDATA = 38'b10110001011110011001100010110111100000;
        11'd372: TDATA = 38'b10110001010010111011111010110111010101;
        11'd373: TDATA = 38'b10110001000111011110110010110111001100;
        11'd374: TDATA = 38'b10110000111100000010011010110111000011;
        11'd375: TDATA = 38'b10110000110000100110100010110110111000;
        11'd376: TDATA = 38'b10110000100101001011010010110110110000;
        11'd377: TDATA = 38'b10110000011001110000100010110110100101;
        11'd378: TDATA = 38'b10110000001110010110100010110110011100;
        11'd379: TDATA = 38'b10110000000010111101000010110110010001;
        11'd380: TDATA = 38'b10101111110111100100001010110110001000;
        11'd381: TDATA = 38'b10101111101100001011111010110110000000;
        11'd382: TDATA = 38'b10101111100000110100010010110101110101;
        11'd383: TDATA = 38'b10101111010101011101010010110101101100;
        11'd384: TDATA = 38'b10101111001010000110110010110101100011;
        11'd385: TDATA = 38'b10101110111110110000111010110101011000;
        11'd386: TDATA = 38'b10101110110011011011101010110101010000;
        11'd387: TDATA = 38'b10101110101000000111000010110101000101;
        11'd388: TDATA = 38'b10101110011100110010111010110100111100;
        11'd389: TDATA = 38'b10101110010001011111011010110100110011;
        11'd390: TDATA = 38'b10101110000110001100100010110100101001;
        11'd391: TDATA = 38'b10101101111010111010010010110100100000;
        11'd392: TDATA = 38'b10101101101111101000100010110100010101;
        11'd393: TDATA = 38'b10101101100100010111011010110100001100;
        11'd394: TDATA = 38'b10101101011001000110111010110100000100;
        11'd395: TDATA = 38'b10101101001101110110111010110011111001;
        11'd396: TDATA = 38'b10101101000010100111101010110011110000;
        11'd397: TDATA = 38'b10101100110111011000111010110011101000;
        11'd398: TDATA = 38'b10101100101100001010101010110011011101;
        11'd399: TDATA = 38'b10101100100000111101001010110011010100;
        11'd400: TDATA = 38'b10101100010101110000001010110011001011;
        11'd401: TDATA = 38'b10101100001010100011110010110011000001;
        11'd402: TDATA = 38'b10101011111111010111111010110010111000;
        11'd403: TDATA = 38'b10101011110100001100101010110010101111;
        11'd404: TDATA = 38'b10101011101001000010000010110010100101;
        11'd405: TDATA = 38'b10101011011101110111111010110010011100;
        11'd406: TDATA = 38'b10101011010010101110011010110010010011;
        11'd407: TDATA = 38'b10101011000111100101100010110010001001;
        11'd408: TDATA = 38'b10101010111100011101001010110010000000;
        11'd409: TDATA = 38'b10101010110001010101100010110001111000;
        11'd410: TDATA = 38'b10101010100110001110010010110001101101;
        11'd411: TDATA = 38'b10101010011011000111101010110001100100;
        11'd412: TDATA = 38'b10101010010000000001101010110001011100;
        11'd413: TDATA = 38'b10101010000100111100010010110001010001;
        11'd414: TDATA = 38'b10101001111001110111011010110001001000;
        11'd415: TDATA = 38'b10101001101110110011001010110001000000;
        11'd416: TDATA = 38'b10101001100011101111011010110000110111;
        11'd417: TDATA = 38'b10101001011000101100010010110000101100;
        11'd418: TDATA = 38'b10101001001101101001101010110000100100;
        11'd419: TDATA = 38'b10101001000010100111110010110000011011;
        11'd420: TDATA = 38'b10101000110111100110010010110000010001;
        11'd421: TDATA = 38'b10101000101100100101011010110000001000;
        11'd422: TDATA = 38'b10101000100001100101001010110000000000;
        11'd423: TDATA = 38'b10101000010110100101100010101111110111;
        11'd424: TDATA = 38'b10101000001011100110011010101111101101;
        11'd425: TDATA = 38'b10101000000000100111110010101111100100;
        11'd426: TDATA = 38'b10100111110101101001110010101111011011;
        11'd427: TDATA = 38'b10100111101010101100011010101111010001;
        11'd428: TDATA = 38'b10100111011111101111100010101111001000;
        11'd429: TDATA = 38'b10100111010100110011001010101111000000;
        11'd430: TDATA = 38'b10100111001001110111011010101110110111;
        11'd431: TDATA = 38'b10100110111110111100010010101110101101;
        11'd432: TDATA = 38'b10100110110100000001101010101110100101;
        11'd433: TDATA = 38'b10100110101001000111101010101110011100;
        11'd434: TDATA = 38'b10100110011110001110001010101110010011;
        11'd435: TDATA = 38'b10100110010011010101010010101110001001;
        11'd436: TDATA = 38'b10100110001000011100111010101110000000;
        11'd437: TDATA = 38'b10100101111101100101000010101101111000;
        11'd438: TDATA = 38'b10100101110010101101111010101101101111;
        11'd439: TDATA = 38'b10100101100111110111001010101101100101;
        11'd440: TDATA = 38'b10100101011101000001000010101101011101;
        11'd441: TDATA = 38'b10100101010010001011100010101101010100;
        11'd442: TDATA = 38'b10100101000111010110100010101101001100;
        11'd443: TDATA = 38'b10100100111100100010000010101101000011;
        11'd444: TDATA = 38'b10100100110001101110001010101100111001;
        11'd445: TDATA = 38'b10100100100110111010110010101100110000;
        11'd446: TDATA = 38'b10100100011100001000000010101100101000;
        11'd447: TDATA = 38'b10100100010001010101110010101100011111;
        11'd448: TDATA = 38'b10100100000110100100001010101100010101;
        11'd449: TDATA = 38'b10100011111011110011000010101100001100;
        11'd450: TDATA = 38'b10100011110001000010011010101100000100;
        11'd451: TDATA = 38'b10100011100110010010011010101011111100;
        11'd452: TDATA = 38'b10100011011011100010111010101011110011;
        11'd453: TDATA = 38'b10100011010000110100000010101011101001;
        11'd454: TDATA = 38'b10100011000110000101101010101011100001;
        11'd455: TDATA = 38'b10100010111011010111110010101011011000;
        11'd456: TDATA = 38'b10100010110000101010100010101011010000;
        11'd457: TDATA = 38'b10100010100101111101110010101011000111;
        11'd458: TDATA = 38'b10100010011011010001101010101010111111;
        11'd459: TDATA = 38'b10100010010000100110000010101010110101;
        11'd460: TDATA = 38'b10100010000101111010111010101010101100;
        11'd461: TDATA = 38'b10100001111011010000011010101010100100;
        11'd462: TDATA = 38'b10100001110000100110011010101010011100;
        11'd463: TDATA = 38'b10100001100101111100111010101010010011;
        11'd464: TDATA = 38'b10100001011011010100000010101010001011;
        11'd465: TDATA = 38'b10100001010000101011101010101010000001;
        11'd466: TDATA = 38'b10100001000110000011110010101001111000;
        11'd467: TDATA = 38'b10100000111011011100100010101001110000;
        11'd468: TDATA = 38'b10100000110000110101110010101001101000;
        11'd469: TDATA = 38'b10100000100110001111100010101001011111;
        11'd470: TDATA = 38'b10100000011011101001111010101001010101;
        11'd471: TDATA = 38'b10100000010001000100110010101001001101;
        11'd472: TDATA = 38'b10100000000110100000001010101001000100;
        11'd473: TDATA = 38'b10011111111011111100000010101000111100;
        11'd474: TDATA = 38'b10011111110001011000100010101000110100;
        11'd475: TDATA = 38'b10011111100110110101100010101000101011;
        11'd476: TDATA = 38'b10011111011100010011001010101000100011;
        11'd477: TDATA = 38'b10011111010001110001001010101000011001;
        11'd478: TDATA = 38'b10011111000111001111110010101000010001;
        11'd479: TDATA = 38'b10011110111100101110111010101000001000;
        11'd480: TDATA = 38'b10011110110010001110101010101000000000;
        11'd481: TDATA = 38'b10011110100111101110110010100111111000;
        11'd482: TDATA = 38'b10011110011101001111100010100111110000;
        11'd483: TDATA = 38'b10011110010010110000110010100111100111;
        11'd484: TDATA = 38'b10011110001000010010101010100111011111;
        11'd485: TDATA = 38'b10011101111101110100111010100111010101;
        11'd486: TDATA = 38'b10011101110011010111110010100111001101;
        11'd487: TDATA = 38'b10011101101000111011001010100111000100;
        11'd488: TDATA = 38'b10011101011110011111001010100110111100;
        11'd489: TDATA = 38'b10011101010100000011100010100110110100;
        11'd490: TDATA = 38'b10011101001001101000100010100110101100;
        11'd491: TDATA = 38'b10011100111111001110000010100110100100;
        11'd492: TDATA = 38'b10011100110100110100000010100110011011;
        11'd493: TDATA = 38'b10011100101010011010100010100110010011;
        11'd494: TDATA = 38'b10011100100000000001101010100110001011;
        11'd495: TDATA = 38'b10011100010101101001010010100110000001;
        11'd496: TDATA = 38'b10011100001011010001010010100101111001;
        11'd497: TDATA = 38'b10011100000000111010000010100101110001;
        11'd498: TDATA = 38'b10011011110110100011001010100101101000;
        11'd499: TDATA = 38'b10011011101100001100110010100101100000;
        11'd500: TDATA = 38'b10011011100001110111000010100101011000;
        11'd501: TDATA = 38'b10011011010111100001101010100101010000;
        11'd502: TDATA = 38'b10011011001101001100111010100101001000;
        11'd503: TDATA = 38'b10011011000010111000101010100101000000;
        11'd504: TDATA = 38'b10011010111000100100111010100100111000;
        11'd505: TDATA = 38'b10011010101110010001110010100100110000;
        11'd506: TDATA = 38'b10011010100011111111000010100100100111;
        11'd507: TDATA = 38'b10011010011001101100111010100100011111;
        11'd508: TDATA = 38'b10011010001111011011001010100100010111;
        11'd509: TDATA = 38'b10011010000101001010000010100100001111;
        11'd510: TDATA = 38'b10011001111010111001011010100100000101;
        11'd511: TDATA = 38'b10011001110000101001010010100011111101;
        11'd512: TDATA = 38'b10011001100110011001101010100011110101;
        11'd513: TDATA = 38'b10011001011100001010100010100011101101;
        11'd514: TDATA = 38'b10011001010001111011111010100011100100;
        11'd515: TDATA = 38'b10011001000111101101111010100011011100;
        11'd516: TDATA = 38'b10011000111101100000010010100011010100;
        11'd517: TDATA = 38'b10011000110011010011010010100011001100;
        11'd518: TDATA = 38'b10011000101001000110101010100011000100;
        11'd519: TDATA = 38'b10011000011110111010101010100010111100;
        11'd520: TDATA = 38'b10011000010100101111000010100010110100;
        11'd521: TDATA = 38'b10011000001010100100000010100010101100;
        11'd522: TDATA = 38'b10011000000000011001100010100010100100;
        11'd523: TDATA = 38'b10010111110110001111100010100010011100;
        11'd524: TDATA = 38'b10010111101100000110000010100010010100;
        11'd525: TDATA = 38'b10010111100001111101000010100010001100;
        11'd526: TDATA = 38'b10010111010111110100100010100010000100;
        11'd527: TDATA = 38'b10010111001101101100100010100001111100;
        11'd528: TDATA = 38'b10010111000011100101000010100001110100;
        11'd529: TDATA = 38'b10010110111001011110000010100001101100;
        11'd530: TDATA = 38'b10010110101111010111100010100001100100;
        11'd531: TDATA = 38'b10010110100101010001100010100001011100;
        11'd532: TDATA = 38'b10010110011011001100000010100001010100;
        11'd533: TDATA = 38'b10010110010001000111000010100001001100;
        11'd534: TDATA = 38'b10010110000111000010100010100001000100;
        11'd535: TDATA = 38'b10010101111100111110100010100000111100;
        11'd536: TDATA = 38'b10010101110010111011000010100000110100;
        11'd537: TDATA = 38'b10010101101000111000000010100000101100;
        11'd538: TDATA = 38'b10010101011110110101100010100000100100;
        11'd539: TDATA = 38'b10010101010100110011100010100000011100;
        11'd540: TDATA = 38'b10010101001010110010000010100000010100;
        11'd541: TDATA = 38'b10010101000000110001000010100000001100;
        11'd542: TDATA = 38'b10010100110110110000100010100000000100;
        11'd543: TDATA = 38'b10010100101100110000100010011111111100;
        11'd544: TDATA = 38'b10010100100010110001000010011111110100;
        11'd545: TDATA = 38'b10010100011000110010000010011111101100;
        11'd546: TDATA = 38'b10010100001110110011011010011111100100;
        11'd547: TDATA = 38'b10010100000100110101011010011111011100;
        11'd548: TDATA = 38'b10010011111010110111111010011111010100;
        11'd549: TDATA = 38'b10010011110000111010110010011111001100;
        11'd550: TDATA = 38'b10010011100110111110001010011111000100;
        11'd551: TDATA = 38'b10010011011101000010001010011110111101;
        11'd552: TDATA = 38'b10010011010011000110100010011110110101;
        11'd553: TDATA = 38'b10010011001001001011011010011110101101;
        11'd554: TDATA = 38'b10010010111111010000110010011110100101;
        11'd555: TDATA = 38'b10010010110101010110101010011110011101;
        11'd556: TDATA = 38'b10010010101011011101000010011110010111;
        11'd557: TDATA = 38'b10010010100001100011111010011110001111;
        11'd558: TDATA = 38'b10010010010111101011001010011110000111;
        11'd559: TDATA = 38'b10010010001101110011000010011101111111;
        11'd560: TDATA = 38'b10010010000011111011010010011101110111;
        11'd561: TDATA = 38'b10010001111010000100001010011101110000;
        11'd562: TDATA = 38'b10010001110000001101011010011101101000;
        11'd563: TDATA = 38'b10010001100110010111001010011101100000;
        11'd564: TDATA = 38'b10010001011100100001011010011101011000;
        11'd565: TDATA = 38'b10010001010010101100000010011101010000;
        11'd566: TDATA = 38'b10010001001000110111010010011101001000;
        11'd567: TDATA = 38'b10010000111111000010111010011101000001;
        11'd568: TDATA = 38'b10010000110101001111001010011100111001;
        11'd569: TDATA = 38'b10010000101011011011110010011100110001;
        11'd570: TDATA = 38'b10010000100001101000111010011100101001;
        11'd571: TDATA = 38'b10010000010111110110011010011100100001;
        11'd572: TDATA = 38'b10010000001110000100100010011100011011;
        11'd573: TDATA = 38'b10010000000100010011000010011100010100;
        11'd574: TDATA = 38'b10001111111010100010001010011100001100;
        11'd575: TDATA = 38'b10001111110000110001101010011100000100;
        11'd576: TDATA = 38'b10001111100111000001100010011011111100;
        11'd577: TDATA = 38'b10001111011101010010000010011011110100;
        11'd578: TDATA = 38'b10001111010011100011000010011011101100;
        11'd579: TDATA = 38'b10001111001001110100011010011011100101;
        11'd580: TDATA = 38'b10001111000000000110010010011011011111;
        11'd581: TDATA = 38'b10001110110110011000101010011011010111;
        11'd582: TDATA = 38'b10001110101100101011011010011011001111;
        11'd583: TDATA = 38'b10001110100010111110110010011011000111;
        11'd584: TDATA = 38'b10001110011001010010100010011011000000;
        11'd585: TDATA = 38'b10001110001111100110110010011010111000;
        11'd586: TDATA = 38'b10001110000101111011011010011010110000;
        11'd587: TDATA = 38'b10001101111100010000101010011010101001;
        11'd588: TDATA = 38'b10001101110010100110010010011010100001;
        11'd589: TDATA = 38'b10001101101000111100011010011010011001;
        11'd590: TDATA = 38'b10001101011111010011000010011010010011;
        11'd591: TDATA = 38'b10001101010101101010000010011010001011;
        11'd592: TDATA = 38'b10001101001100000001100010011010000100;
        11'd593: TDATA = 38'b10001101000010011001100010011001111100;
        11'd594: TDATA = 38'b10001100111000110010000010011001110100;
        11'd595: TDATA = 38'b10001100101111001010111010011001101101;
        11'd596: TDATA = 38'b10001100100101100100010010011001100101;
        11'd597: TDATA = 38'b10001100011011111110001010011001011101;
        11'd598: TDATA = 38'b10001100010010011000100010011001010111;
        11'd599: TDATA = 38'b10001100001000110011010010011001010000;
        11'd600: TDATA = 38'b10001011111111001110100010011001001000;
        11'd601: TDATA = 38'b10001011110101101010010010011001000000;
        11'd602: TDATA = 38'b10001011101100000110011010011000111001;
        11'd603: TDATA = 38'b10001011100010100011000010011000110001;
        11'd604: TDATA = 38'b10001011011001000000001010011000101011;
        11'd605: TDATA = 38'b10001011001111011101101010011000100100;
        11'd606: TDATA = 38'b10001011000101111011101010011000011100;
        11'd607: TDATA = 38'b10001010111100011010001010011000010100;
        11'd608: TDATA = 38'b10001010110010111001000010011000001100;
        11'd609: TDATA = 38'b10001010101001011000100010011000000101;
        11'd610: TDATA = 38'b10001010011111111000010010010111111111;
        11'd611: TDATA = 38'b10001010010110011000101010010111111000;
        11'd612: TDATA = 38'b10001010001100111001011010010111110000;
        11'd613: TDATA = 38'b10001010000011011010101010010111101000;
        11'd614: TDATA = 38'b10001001111001111100010010010111100000;
        11'd615: TDATA = 38'b10001001110000011110011010010111011001;
        11'd616: TDATA = 38'b10001001100111000001000010010111010100;
        11'd617: TDATA = 38'b10001001011101100100000010010111001100;
        11'd618: TDATA = 38'b10001001010100000111100010010111000100;
        11'd619: TDATA = 38'b10001001001010101011011010010110111100;
        11'd620: TDATA = 38'b10001001000001001111111010010110110101;
        11'd621: TDATA = 38'b10001000110111110100101010010110101111;
        11'd622: TDATA = 38'b10001000101110011010000010010110101000;
        11'd623: TDATA = 38'b10001000100100111111110010010110100000;
        11'd624: TDATA = 38'b10001000011011100110000010010110011000;
        11'd625: TDATA = 38'b10001000010010001100101010010110010001;
        11'd626: TDATA = 38'b10001000001000110011110010010110001011;
        11'd627: TDATA = 38'b10000111111111011011010010010110000100;
        11'd628: TDATA = 38'b10000111110110000011010010010101111100;
        11'd629: TDATA = 38'b10000111101100101011110010010101110100;
        11'd630: TDATA = 38'b10000111100011010100101010010101101101;
        11'd631: TDATA = 38'b10000111011001111110000010010101100111;
        11'd632: TDATA = 38'b10000111010000100111110010010101100000;
        11'd633: TDATA = 38'b10000111000111010010000010010101011000;
        11'd634: TDATA = 38'b10000110111101111100101010010101010000;
        11'd635: TDATA = 38'b10000110110100100111110010010101001001;
        11'd636: TDATA = 38'b10000110101011010011011010010101000100;
        11'd637: TDATA = 38'b10000110100001111111011010010100111100;
        11'd638: TDATA = 38'b10000110011000101011111010010100110100;
        11'd639: TDATA = 38'b10000110001111011000110010010100101101;
        11'd640: TDATA = 38'b10000110000110000110001010010100100111;
        11'd641: TDATA = 38'b10000101111100110011111010010100100000;
        11'd642: TDATA = 38'b10000101110011100010001010010100011000;
        11'd643: TDATA = 38'b10000101101010010000110010010100010001;
        11'd644: TDATA = 38'b10000101100000111111111010010100001001;
        11'd645: TDATA = 38'b10000101010111101111100010010100000100;
        11'd646: TDATA = 38'b10000101001110011111100010010011111100;
        11'd647: TDATA = 38'b10000101000101001111111010010011110101;
        11'd648: TDATA = 38'b10000100111100000000110010010011101111;
        11'd649: TDATA = 38'b10000100110010110010001010010011100111;
        11'd650: TDATA = 38'b10000100101001100011111010010011100000;
        11'd651: TDATA = 38'b10000100100000010110000010010011011001;
        11'd652: TDATA = 38'b10000100010111001000101010010011010011;
        11'd653: TDATA = 38'b10000100001101111011110010010011001011;
        11'd654: TDATA = 38'b10000100000100101111001010010011000100;
        11'd655: TDATA = 38'b10000011111011100011001010010010111101;
        11'd656: TDATA = 38'b10000011110010010111100010010010110111;
        11'd657: TDATA = 38'b10000011101001001100010010010010110000;
        11'd658: TDATA = 38'b10000011100000000001100010010010101000;
        11'd659: TDATA = 38'b10000011010110110111001010010010100001;
        11'd660: TDATA = 38'b10000011001101101101010010010010011011;
        11'd661: TDATA = 38'b10000011000100100011111010010010010100;
        11'd662: TDATA = 38'b10000010111011011010110010010010001100;
        11'd663: TDATA = 38'b10000010110010010010001010010010000101;
        11'd664: TDATA = 38'b10000010101001001010000010010010000000;
        11'd665: TDATA = 38'b10000010100000000010010010010001111000;
        11'd666: TDATA = 38'b10000010010110111011000010010001110000;
        11'd667: TDATA = 38'b10000010001101110100001010010001101011;
        11'd668: TDATA = 38'b10000010000100101101101010010001100100;
        11'd669: TDATA = 38'b10000001111011100111101010010001011100;
        11'd670: TDATA = 38'b10000001110010100010000010010001010101;
        11'd671: TDATA = 38'b10000001101001011100111010010001001111;
        11'd672: TDATA = 38'b10000001100000011000001010010001001000;
        11'd673: TDATA = 38'b10000001010111010011110010010001000001;
        11'd674: TDATA = 38'b10000001001110001111111010010000111011;
        11'd675: TDATA = 38'b10000001000101001100011010010000110100;
        11'd676: TDATA = 38'b10000000111100001001011010010000101101;
        11'd677: TDATA = 38'b10000000110011000110110010010000100111;
        11'd678: TDATA = 38'b10000000101010000100101010010000100000;
        11'd679: TDATA = 38'b10000000100001000010111010010000011000;
        11'd680: TDATA = 38'b10000000011000000001100010010000010011;
        11'd681: TDATA = 38'b10000000001111000000101010010000001100;
        11'd682: TDATA = 38'b10000000000110000000001010010000000100;
        11'd683: TDATA = 38'b01111111111101000000000010001111111101;
        11'd684: TDATA = 38'b01111111110100000000011010001111111000;
        11'd685: TDATA = 38'b01111111101011000001001010001111110000;
        11'd686: TDATA = 38'b01111111100010000010011010001111101001;
        11'd687: TDATA = 38'b01111111011001000100000010001111100011;
        11'd688: TDATA = 38'b01111111010000000110000010001111011100;
        11'd689: TDATA = 38'b01111111000111001000100010001111010101;
        11'd690: TDATA = 38'b01111110111110001011011010001111001111;
        11'd691: TDATA = 38'b01111110110101001110101010001111001000;
        11'd692: TDATA = 38'b01111110101100010010010010001111000001;
        11'd693: TDATA = 38'b01111110100011010110100010001110111011;
        11'd694: TDATA = 38'b01111110011010011011000010001110110100;
        11'd695: TDATA = 38'b01111110010001100000000010001110101100;
        11'd696: TDATA = 38'b01111110001000100101011010001110100111;
        11'd697: TDATA = 38'b01111101111111101011001010001110100000;
        11'd698: TDATA = 38'b01111101110110110001011010001110011000;
        11'd699: TDATA = 38'b01111101101101111000000010001110010011;
        11'd700: TDATA = 38'b01111101100100111111000010001110001100;
        11'd701: TDATA = 38'b01111101011100000110011010001110000101;
        11'd702: TDATA = 38'b01111101010011001110010010001101111111;
        11'd703: TDATA = 38'b01111101001010010110101010001101111000;
        11'd704: TDATA = 38'b01111101000001011111010010001101110001;
        11'd705: TDATA = 38'b01111100111000101000011010001101101011;
        11'd706: TDATA = 38'b01111100101111110001111010001101100100;
        11'd707: TDATA = 38'b01111100100110111011110010001101011101;
        11'd708: TDATA = 38'b01111100011110000110001010001101011000;
        11'd709: TDATA = 38'b01111100010101010000111010001101010000;
        11'd710: TDATA = 38'b01111100001100011100000010001101001001;
        11'd711: TDATA = 38'b01111100000011100111101010001101000100;
        11'd712: TDATA = 38'b01111011111010110011101010001100111100;
        11'd713: TDATA = 38'b01111011110010000000000010001100110111;
        11'd714: TDATA = 38'b01111011101001001100110010001100110000;
        11'd715: TDATA = 38'b01111011100000011010000010001100101001;
        11'd716: TDATA = 38'b01111011010111100111100010001100100011;
        11'd717: TDATA = 38'b01111011001110110101100010001100011100;
        11'd718: TDATA = 38'b01111011000110000100000010001100010111;
        11'd719: TDATA = 38'b01111010111101010010110010001100010000;
        11'd720: TDATA = 38'b01111010110100100010000010001100001000;
        11'd721: TDATA = 38'b01111010101011110001101010001100000011;
        11'd722: TDATA = 38'b01111010100011000001110010001011111100;
        11'd723: TDATA = 38'b01111010011010010010001010001011110101;
        11'd724: TDATA = 38'b01111010010001100011000010001011101111;
        11'd725: TDATA = 38'b01111010001000110100010010001011101000;
        11'd726: TDATA = 38'b01111010000000000101111010001011100011;
        11'd727: TDATA = 38'b01111001110111011000000010001011011100;
        11'd728: TDATA = 38'b01111001101110101010011010001011010100;
        11'd729: TDATA = 38'b01111001100101111101010010001011001111;
        11'd730: TDATA = 38'b01111001011101010000100010001011001000;
        11'd731: TDATA = 38'b01111001010100100100010010001011000001;
        11'd732: TDATA = 38'b01111001001011111000010010001010111100;
        11'd733: TDATA = 38'b01111001000011001100110010001010110101;
        11'd734: TDATA = 38'b01111000111010100001101010001010101111;
        11'd735: TDATA = 38'b01111000110001110110111010001010101000;
        11'd736: TDATA = 38'b01111000101001001100100010001010100011;
        11'd737: TDATA = 38'b01111000100000100010100010001010011100;
        11'd738: TDATA = 38'b01111000010111111001000010001010010100;
        11'd739: TDATA = 38'b01111000001111001111111010001010010000;
        11'd740: TDATA = 38'b01111000000110100111001010001010001000;
        11'd741: TDATA = 38'b01110111111101111110110010001010000001;
        11'd742: TDATA = 38'b01110111110101010110110010001001111100;
        11'd743: TDATA = 38'b01110111101100101111010010001001110101;
        11'd744: TDATA = 38'b01110111100100001000001010001001110000;
        11'd745: TDATA = 38'b01110111011011100001010010001001101000;
        11'd746: TDATA = 38'b01110111010010111010111010001001100011;
        11'd747: TDATA = 38'b01110111001010010100111010001001011100;
        11'd748: TDATA = 38'b01110111000001101111011010001001010101;
        11'd749: TDATA = 38'b01110110111001001010001010001001010000;
        11'd750: TDATA = 38'b01110110110000100101011010001001001001;
        11'd751: TDATA = 38'b01110110101000000000111010001001000100;
        11'd752: TDATA = 38'b01110110011111011100111010001000111100;
        11'd753: TDATA = 38'b01110110010110111001010010001000110111;
        11'd754: TDATA = 38'b01110110001110010110000010001000110000;
        11'd755: TDATA = 38'b01110110000101110011001010001000101001;
        11'd756: TDATA = 38'b01110101111101010000110010001000100100;
        11'd757: TDATA = 38'b01110101110100101110101010001000011101;
        11'd758: TDATA = 38'b01110101101100001101000010001000011000;
        11'd759: TDATA = 38'b01110101100011101011101010001000010001;
        11'd760: TDATA = 38'b01110101011011001010110010001000001100;
        11'd761: TDATA = 38'b01110101010010101010010010001000000100;
        11'd762: TDATA = 38'b01110101001010001010001010000111111111;
        11'd763: TDATA = 38'b01110101000001101010011010000111111000;
        11'd764: TDATA = 38'b01110100111001001011000010000111110011;
        11'd765: TDATA = 38'b01110100110000101100000010000111101100;
        11'd766: TDATA = 38'b01110100101000001101100010000111100111;
        11'd767: TDATA = 38'b01110100011111101111010010000111100000;
        11'd768: TDATA = 38'b01110100010111010001100010000111011001;
        11'd769: TDATA = 38'b01110100001110110100000010000111010100;
        11'd770: TDATA = 38'b01110100000110010111000010000111001101;
        11'd771: TDATA = 38'b01110011111101111010011010000111000111;
        11'd772: TDATA = 38'b01110011110101011110000010000111000001;
        11'd773: TDATA = 38'b01110011101101000010001010000110111100;
        11'd774: TDATA = 38'b01110011100100100110101010000110110100;
        11'd775: TDATA = 38'b01110011011100001011100010000110101111;
        11'd776: TDATA = 38'b01110011010011110000110010000110101000;
        11'd777: TDATA = 38'b01110011001011010110011010000110100011;
        11'd778: TDATA = 38'b01110011000010111100011010000110011100;
        11'd779: TDATA = 38'b01110010111010100010111010000110010111;
        11'd780: TDATA = 38'b01110010110010001001101010000110010000;
        11'd781: TDATA = 38'b01110010101001110000110010000110001001;
        11'd782: TDATA = 38'b01110010100001011000010010000110000100;
        11'd783: TDATA = 38'b01110010011001000000010010000101111111;
        11'd784: TDATA = 38'b01110010010000101000100010000101111000;
        11'd785: TDATA = 38'b01110010001000010001001010000101110011;
        11'd786: TDATA = 38'b01110001111111111010010010000101101100;
        11'd787: TDATA = 38'b01110001110111100011101010000101100101;
        11'd788: TDATA = 38'b01110001101111001101100010000101100000;
        11'd789: TDATA = 38'b01110001100110110111101010000101011001;
        11'd790: TDATA = 38'b01110001011110100010001010000101010100;
        11'd791: TDATA = 38'b01110001010110001101001010000101001101;
        11'd792: TDATA = 38'b01110001001101111000011010000101001000;
        11'd793: TDATA = 38'b01110001000101100100001010000101000001;
        11'd794: TDATA = 38'b01110000111101010000001010000100111100;
        11'd795: TDATA = 38'b01110000110100111100101010000100110101;
        11'd796: TDATA = 38'b01110000101100101001011010000100110000;
        11'd797: TDATA = 38'b01110000100100010110101010000100101001;
        11'd798: TDATA = 38'b01110000011100000100001010000100100100;
        11'd799: TDATA = 38'b01110000010011110010001010000100011101;
        11'd800: TDATA = 38'b01110000001011100000011010000100011000;
        11'd801: TDATA = 38'b01110000000011001111000010000100010011;
        11'd802: TDATA = 38'b01101111111010111110001010000100001100;
        11'd803: TDATA = 38'b01101111110010101101100010000100000101;
        11'd804: TDATA = 38'b01101111101010011101010010000100000000;
        11'd805: TDATA = 38'b01101111100010001101011010000011111011;
        11'd806: TDATA = 38'b01101111011001111101111010000011110100;
        11'd807: TDATA = 38'b01101111010001101110111010000011101111;
        11'd808: TDATA = 38'b01101111001001100000001010000011101000;
        11'd809: TDATA = 38'b01101111000001010001110010000011100011;
        11'd810: TDATA = 38'b01101110111001000011110010000011011101;
        11'd811: TDATA = 38'b01101110110000110110001010000011010111;
        11'd812: TDATA = 38'b01101110101000101000111010000011010000;
        11'd813: TDATA = 38'b01101110100000011011111010000011001100;
        11'd814: TDATA = 38'b01101110011000001111011010000011000101;
        11'd815: TDATA = 38'b01101110010000000011010010000011000000;
        11'd816: TDATA = 38'b01101110000111110111011010000010111001;
        11'd817: TDATA = 38'b01101101111111101100000010000010110100;
        11'd818: TDATA = 38'b01101101110111100000111010000010101101;
        11'd819: TDATA = 38'b01101101101111010110010010000010101000;
        11'd820: TDATA = 38'b01101101100111001011111010000010100011;
        11'd821: TDATA = 38'b01101101011111000001111010000010011100;
        11'd822: TDATA = 38'b01101101010110111000010010000010010111;
        11'd823: TDATA = 38'b01101101001110101111000010000010010000;
        11'd824: TDATA = 38'b01101101000110100110001010000010001011;
        11'd825: TDATA = 38'b01101100111110011101101010000010000101;
        11'd826: TDATA = 38'b01101100110110010101100010000010000000;
        11'd827: TDATA = 38'b01101100101110001101101010000001111001;
        11'd828: TDATA = 38'b01101100100110000110010010000001110100;
        11'd829: TDATA = 38'b01101100011101111111001010000001101101;
        11'd830: TDATA = 38'b01101100010101111000100010000001101000;
        11'd831: TDATA = 38'b01101100001101110010001010000001100011;
        11'd832: TDATA = 38'b01101100000101101100001010000001011100;
        11'd833: TDATA = 38'b01101011111101100110100010000001010111;
        11'd834: TDATA = 38'b01101011110101100001001010000001010001;
        11'd835: TDATA = 38'b01101011101101011100010010000001001100;
        11'd836: TDATA = 38'b01101011100101010111110010000001000101;
        11'd837: TDATA = 38'b01101011011101010011100010000001000000;
        11'd838: TDATA = 38'b01101011010101001111101010000000111011;
        11'd839: TDATA = 38'b01101011001101001100001010000000110100;
        11'd840: TDATA = 38'b01101011000101001001000010000000110000;
        11'd841: TDATA = 38'b01101010111101000110010010000000101001;
        11'd842: TDATA = 38'b01101010110101000011111010000000100100;
        11'd843: TDATA = 38'b01101010101101000001110010000000011111;
        11'd844: TDATA = 38'b01101010100101000000001010000000011000;
        11'd845: TDATA = 38'b01101010011100111110110010000000010011;
        11'd846: TDATA = 38'b01101010010100111101110010000000001100;
        11'd847: TDATA = 38'b01101010001100111101001010000000000111;
        11'd848: TDATA = 38'b01101010000100111100111010000000000001;
        11'd849: TDATA = 38'b01101001111100111100111001111111111100;
        11'd850: TDATA = 38'b01101001110100111101010001111111110101;
        11'd851: TDATA = 38'b01101001101100111110001001111111110000;
        11'd852: TDATA = 38'b01101001100100111111010001111111101011;
        11'd853: TDATA = 38'b01101001011101000000101001111111100101;
        11'd854: TDATA = 38'b01101001010101000010100001111111100000;
        11'd855: TDATA = 38'b01101001001101000100110001111111011011;
        11'd856: TDATA = 38'b01101001000101000111010001111111010100;
        11'd857: TDATA = 38'b01101000111101001010001001111111001111;
        11'd858: TDATA = 38'b01101000110101001101011001111111001001;
        11'd859: TDATA = 38'b01101000101101010000111001111111000100;
        11'd860: TDATA = 38'b01101000100101010100111001111110111111;
        11'd861: TDATA = 38'b01101000011101011001001001111110111000;
        11'd862: TDATA = 38'b01101000010101011101110001111110110011;
        11'd863: TDATA = 38'b01101000001101100010110001111110101101;
        11'd864: TDATA = 38'b01101000000101101000001001111110101000;
        11'd865: TDATA = 38'b01100111111101101101110001111110100001;
        11'd866: TDATA = 38'b01100111110101110011110001111110011100;
        11'd867: TDATA = 38'b01100111101101111010001001111110010111;
        11'd868: TDATA = 38'b01100111100110000000111001111110010001;
        11'd869: TDATA = 38'b01100111011110001000000001111110001100;
        11'd870: TDATA = 38'b01100111010110001111011001111110000111;
        11'd871: TDATA = 38'b01100111001110010111001001111110000000;
        11'd872: TDATA = 38'b01100111000110011111010001111101111100;
        11'd873: TDATA = 38'b01100110111110100111101001111101110101;
        11'd874: TDATA = 38'b01100110110110110000100001111101110000;
        11'd875: TDATA = 38'b01100110101110111001101001111101101011;
        11'd876: TDATA = 38'b01100110100111000011001001111101100101;
        11'd877: TDATA = 38'b01100110011111001100111001111101100000;
        11'd878: TDATA = 38'b01100110010111010111000001111101011011;
        11'd879: TDATA = 38'b01100110001111100001101001111101010100;
        11'd880: TDATA = 38'b01100110000111101100011001111101010000;
        11'd881: TDATA = 38'b01100101111111110111101001111101001001;
        11'd882: TDATA = 38'b01100101111000000011001001111101000100;
        11'd883: TDATA = 38'b01100101110000001111000001111101000000;
        11'd884: TDATA = 38'b01100101101000011011010001111100111001;
        11'd885: TDATA = 38'b01100101100000100111110001111100110100;
        11'd886: TDATA = 38'b01100101011000110100110001111100101111;
        11'd887: TDATA = 38'b01100101010001000010000001111100101001;
        11'd888: TDATA = 38'b01100101001001001111100001111100100100;
        11'd889: TDATA = 38'b01100101000001011101100001111100011111;
        11'd890: TDATA = 38'b01100100111001101011110001111100011000;
        11'd891: TDATA = 38'b01100100110001111010010001111100010100;
        11'd892: TDATA = 38'b01100100101010001001010001111100001111;
        11'd893: TDATA = 38'b01100100100010011000100001111100001000;
        11'd894: TDATA = 38'b01100100011010101000001001111100000100;
        11'd895: TDATA = 38'b01100100010010111000001001111011111101;
        11'd896: TDATA = 38'b01100100001011001000011001111011111000;
        11'd897: TDATA = 38'b01100100000011011001000001111011110100;
        11'd898: TDATA = 38'b01100011111011101001111001111011101101;
        11'd899: TDATA = 38'b01100011110011111011010001111011101000;
        11'd900: TDATA = 38'b01100011101100001100111001111011100100;
        11'd901: TDATA = 38'b01100011100100011110111001111011011101;
        11'd902: TDATA = 38'b01100011011100110001001001111011011000;
        11'd903: TDATA = 38'b01100011010101000011110001111011010100;
        11'd904: TDATA = 38'b01100011001101010110110001111011001101;
        11'd905: TDATA = 38'b01100011000101101010000001111011001000;
        11'd906: TDATA = 38'b01100010111101111101101001111011000011;
        11'd907: TDATA = 38'b01100010110110010001101001111010111101;
        11'd908: TDATA = 38'b01100010101110100101111001111010111000;
        11'd909: TDATA = 38'b01100010100110111010101001111010110011;
        11'd910: TDATA = 38'b01100010011111001111100001111010101101;
        11'd911: TDATA = 38'b01100010010111100100111001111010101000;
        11'd912: TDATA = 38'b01100010001111111010100001111010100011;
        11'd913: TDATA = 38'b01100010001000010000011001111010011101;
        11'd914: TDATA = 38'b01100010000000100110110001111010011000;
        11'd915: TDATA = 38'b01100001111000111101011001111010010011;
        11'd916: TDATA = 38'b01100001110001010100010001111010001101;
        11'd917: TDATA = 38'b01100001101001101011101001111010001000;
        11'd918: TDATA = 38'b01100001100010000011010001111010000100;
        11'd919: TDATA = 38'b01100001011010011011001001111001111101;
        11'd920: TDATA = 38'b01100001010010110011011001111001111000;
        11'd921: TDATA = 38'b01100001001011001100000001111001110100;
        11'd922: TDATA = 38'b01100001000011100100111001111001101111;
        11'd923: TDATA = 38'b01100000111011111110010001111001101000;
        11'd924: TDATA = 38'b01100000110100010111110001111001100100;
        11'd925: TDATA = 38'b01100000101100110001101001111001011111;
        11'd926: TDATA = 38'b01100000100101001011111001111001011001;
        11'd927: TDATA = 38'b01100000011101100110100001111001010100;
        11'd928: TDATA = 38'b01100000010110000001011001111001010000;
        11'd929: TDATA = 38'b01100000001110011100101001111001001001;
        11'd930: TDATA = 38'b01100000000110111000001001111001000100;
        11'd931: TDATA = 38'b01011111111111010100000001111001000000;
        11'd932: TDATA = 38'b01011111110111110000010001111000111001;
        11'd933: TDATA = 38'b01011111110000001100110001111000110101;
        11'd934: TDATA = 38'b01011111101000101001100001111000110000;
        11'd935: TDATA = 38'b01011111100001000110110001111000101011;
        11'd936: TDATA = 38'b01011111011001100100010001111000100101;
        11'd937: TDATA = 38'b01011111010010000010000001111000100000;
        11'd938: TDATA = 38'b01011111001010100000001001111000011011;
        11'd939: TDATA = 38'b01011111000010111110101001111000010101;
        11'd940: TDATA = 38'b01011110111011011101011001111000010000;
        11'd941: TDATA = 38'b01011110110011111100100001111000001100;
        11'd942: TDATA = 38'b01011110101100011011111001111000000111;
        11'd943: TDATA = 38'b01011110100100111011101001111000000000;
        11'd944: TDATA = 38'b01011110011101011011110001110111111100;
        11'd945: TDATA = 38'b01011110010101111100001001110111110111;
        11'd946: TDATA = 38'b01011110001110011100111001110111110001;
        11'd947: TDATA = 38'b01011110000110111101111001110111101100;
        11'd948: TDATA = 38'b01011101111111011111010001110111101000;
        11'd949: TDATA = 38'b01011101111000000000111001110111100011;
        11'd950: TDATA = 38'b01011101110000100010111001110111011101;
        11'd951: TDATA = 38'b01011101101001000101001001110111011000;
        11'd952: TDATA = 38'b01011101100001100111110001110111010100;
        11'd953: TDATA = 38'b01011101011010001010110001110111001111;
        11'd954: TDATA = 38'b01011101010010101110000001110111001000;
        11'd955: TDATA = 38'b01011101001011010001100001110111000100;
        11'd956: TDATA = 38'b01011101000011110101011001110110111111;
        11'd957: TDATA = 38'b01011100111100011001101001110110111001;
        11'd958: TDATA = 38'b01011100110100111110001001110110110100;
        11'd959: TDATA = 38'b01011100101101100011000001110110110000;
        11'd960: TDATA = 38'b01011100100110001000001001110110101011;
        11'd961: TDATA = 38'b01011100011110101101101001110110100101;
        11'd962: TDATA = 38'b01011100010111010011011001110110100000;
        11'd963: TDATA = 38'b01011100001111111001100001110110011100;
        11'd964: TDATA = 38'b01011100001000100000000001110110010111;
        11'd965: TDATA = 38'b01011100000001000110110001110110010001;
        11'd966: TDATA = 38'b01011011111001101101110001110110001100;
        11'd967: TDATA = 38'b01011011110010010101001001110110001000;
        11'd968: TDATA = 38'b01011011101010111100110001110110000011;
        11'd969: TDATA = 38'b01011011100011100100110001110101111101;
        11'd970: TDATA = 38'b01011011011100001101001001110101111000;
        11'd971: TDATA = 38'b01011011010100110101101001110101110100;
        11'd972: TDATA = 38'b01011011001101011110101001110101101111;
        11'd973: TDATA = 38'b01011011000110000111111001110101101001;
        11'd974: TDATA = 38'b01011010111110110001011001110101100100;
        11'd975: TDATA = 38'b01011010110111011011010001110101100000;
        11'd976: TDATA = 38'b01011010110000000101011001110101011011;
        11'd977: TDATA = 38'b01011010101000101111111001110101010101;
        11'd978: TDATA = 38'b01011010100001011010110001110101010000;
        11'd979: TDATA = 38'b01011010011010000101110001110101001100;
        11'd980: TDATA = 38'b01011010010010110001010001110101000111;
        11'd981: TDATA = 38'b01011010001011011100111001110101000001;
        11'd982: TDATA = 38'b01011010000100001001000001110100111100;
        11'd983: TDATA = 38'b01011001111100110101010001110100111000;
        11'd984: TDATA = 38'b01011001110101100010000001110100110011;
        11'd985: TDATA = 38'b01011001101110001110111001110100101111;
        11'd986: TDATA = 38'b01011001100110111100001001110100101000;
        11'd987: TDATA = 38'b01011001011111101001110001110100100100;
        11'd988: TDATA = 38'b01011001011000010111101001110100100000;
        11'd989: TDATA = 38'b01011001010001000101110001110100011011;
        11'd990: TDATA = 38'b01011001001001110100010001110100010101;
        11'd991: TDATA = 38'b01011001000010100011001001110100010000;
        11'd992: TDATA = 38'b01011000111011010010010001110100001100;
        11'd993: TDATA = 38'b01011000110100000001101001110100000111;
        11'd994: TDATA = 38'b01011000101100110001011001110100000001;
        11'd995: TDATA = 38'b01011000100101100001011001110011111100;
        11'd996: TDATA = 38'b01011000011110010001101001110011111000;
        11'd997: TDATA = 38'b01011000010111000010010001110011110100;
        11'd998: TDATA = 38'b01011000001111110011010001110011101111;
        11'd999: TDATA = 38'b01011000001000100100100001110011101001;
        11'd1000: TDATA = 38'b01011000000001010110000001110011100100;
        11'd1001: TDATA = 38'b01010111111010000111111001110011100000;
        11'd1002: TDATA = 38'b01010111110010111010000001110011011011;
        11'd1003: TDATA = 38'b01010111101011101100100001110011010101;
        11'd1004: TDATA = 38'b01010111100100011111010001110011010001;
        11'd1005: TDATA = 38'b01010111011101010010010001110011001100;
        11'd1006: TDATA = 38'b01010111010110000101101001110011001000;
        11'd1007: TDATA = 38'b01010111001110111001010001110011000011;
        11'd1008: TDATA = 38'b01010111000111101101010001110010111101;
        11'd1009: TDATA = 38'b01010111000000100001100001110010111001;
        11'd1010: TDATA = 38'b01010110111001010110000001110010110100;
        11'd1011: TDATA = 38'b01010110110010001010111001110010110000;
        11'd1012: TDATA = 38'b01010110101011000000001001110010101100;
        11'd1013: TDATA = 38'b01010110100011110101100001110010100101;
        11'd1014: TDATA = 38'b01010110011100101011010001110010100000;
        11'd1015: TDATA = 38'b01010110010101100001011001110010011100;
        11'd1016: TDATA = 38'b01010110001110010111110001110010011000;
        11'd1017: TDATA = 38'b01010110000111001110011001110010010011;
        11'd1018: TDATA = 38'b01010110000000000101011001110010001111;
        11'd1019: TDATA = 38'b01010101111000111100101001110010001000;
        11'd1020: TDATA = 38'b01010101110001110100001001110010000100;
        11'd1021: TDATA = 38'b01010101101010101100000001110010000000;
        11'd1022: TDATA = 38'b01010101100011100100001001110001111011;
        11'd1023: TDATA = 38'b01010101011100011100101001110001110111;
        11'd1024: TDATA = 38'b01010101010101010101011001110001110001;
        11'd1025: TDATA = 38'b01010101001110001110011001110001101100;
        11'd1026: TDATA = 38'b01010101000111000111110001110001101000;
        11'd1027: TDATA = 38'b01010101000000000001011001110001100100;
        11'd1028: TDATA = 38'b01010100111000111011010001110001011111;
        11'd1029: TDATA = 38'b01010100110001110101100001110001011001;
        11'd1030: TDATA = 38'b01010100101010110000000001110001010100;
        11'd1031: TDATA = 38'b01010100100011101010110001110001010000;
        11'd1032: TDATA = 38'b01010100011100100101111001110001001100;
        11'd1033: TDATA = 38'b01010100010101100001010001110001000111;
        11'd1034: TDATA = 38'b01010100001110011101000001110001000011;
        11'd1035: TDATA = 38'b01010100000111011001000001110000111101;
        11'd1036: TDATA = 38'b01010100000000010101010001110000111001;
        11'd1037: TDATA = 38'b01010011111001010001111001110000110100;
        11'd1038: TDATA = 38'b01010011110010001110101001110000110000;
        11'd1039: TDATA = 38'b01010011101011001011111001110000101100;
        11'd1040: TDATA = 38'b01010011100100001001010001110000100111;
        11'd1041: TDATA = 38'b01010011011101000111000001110000100001;
        11'd1042: TDATA = 38'b01010011010110000101000001110000011101;
        11'd1043: TDATA = 38'b01010011001111000011011001110000011000;
        11'd1044: TDATA = 38'b01010011001000000010000001110000010100;
        11'd1045: TDATA = 38'b01010011000001000000111001110000010000;
        11'd1046: TDATA = 38'b01010010111010000000001001110000001011;
        11'd1047: TDATA = 38'b01010010110010111111101001110000000101;
        11'd1048: TDATA = 38'b01010010101011111111011001110000000000;
        11'd1049: TDATA = 38'b01010010100100111111011001101111111100;
        11'd1050: TDATA = 38'b01010010011101111111110001101111111000;
        11'd1051: TDATA = 38'b01010010010111000000011001101111110100;
        11'd1052: TDATA = 38'b01010010010000000001011001101111101111;
        11'd1053: TDATA = 38'b01010010001001000010100001101111101011;
        11'd1054: TDATA = 38'b01010010000010000100000001101111100101;
        11'd1055: TDATA = 38'b01010001111011000101111001101111100000;
        11'd1056: TDATA = 38'b01010001110100000111111001101111011100;
        11'd1057: TDATA = 38'b01010001101101001010010001101111011000;
        11'd1058: TDATA = 38'b01010001100110001101000001101111010100;
        11'd1059: TDATA = 38'b01010001011111001111111001101111001111;
        11'd1060: TDATA = 38'b01010001011000010011001001101111001001;
        11'd1061: TDATA = 38'b01010001010001010110101001101111000101;
        11'd1062: TDATA = 38'b01010001001010011010011001101111000000;
        11'd1063: TDATA = 38'b01010001000011011110100001101110111100;
        11'd1064: TDATA = 38'b01010000111100100010111001101110111000;
        11'd1065: TDATA = 38'b01010000110101100111100001101110110011;
        11'd1066: TDATA = 38'b01010000101110101100100001101110101111;
        11'd1067: TDATA = 38'b01010000100111110001110001101110101001;
        11'd1068: TDATA = 38'b01010000100000110111010001101110100101;
        11'd1069: TDATA = 38'b01010000011001111101000001101110100000;
        11'd1070: TDATA = 38'b01010000010011000011001001101110011100;
        11'd1071: TDATA = 38'b01010000001100001001100001101110011000;
        11'd1072: TDATA = 38'b01010000000101010000001001101110010100;
        11'd1073: TDATA = 38'b01001111111110010111000001101110001111;
        11'd1074: TDATA = 38'b01001111110111011110010001101110001011;
        11'd1075: TDATA = 38'b01001111110000100101110001101110000101;
        11'd1076: TDATA = 38'b01001111101001101101100001101110000000;
        11'd1077: TDATA = 38'b01001111100010110101100001101101111100;
        11'd1078: TDATA = 38'b01001111011011111101111001101101111000;
        11'd1079: TDATA = 38'b01001111010101000110100001101101110100;
        11'd1080: TDATA = 38'b01001111001110001111011001101101110000;
        11'd1081: TDATA = 38'b01001111000111011000101001101101101011;
        11'd1082: TDATA = 38'b01001111000000100010000001101101100111;
        11'd1083: TDATA = 38'b01001110111001101011110001101101100001;
        11'd1084: TDATA = 38'b01001110110010110101110001101101011100;
        11'd1085: TDATA = 38'b01001110101100000000001001101101011000;
        11'd1086: TDATA = 38'b01001110100101001010101001101101010100;
        11'd1087: TDATA = 38'b01001110011110010101100001101101010000;
        11'd1088: TDATA = 38'b01001110010111100000101001101101001100;
        11'd1089: TDATA = 38'b01001110010000101100001001101101000111;
        11'd1090: TDATA = 38'b01001110001001110111110001101101000011;
        11'd1091: TDATA = 38'b01001110000011000011110001101100111111;
        11'd1092: TDATA = 38'b01001101111100010000000001101100111001;
        11'd1093: TDATA = 38'b01001101110101011100100001101100110101;
        11'd1094: TDATA = 38'b01001101101110101001010001101100110000;
        11'd1095: TDATA = 38'b01001101100111110110011001101100101100;
        11'd1096: TDATA = 38'b01001101100001000011110001101100101000;
        11'd1097: TDATA = 38'b01001101011010010001011001101100100100;
        11'd1098: TDATA = 38'b01001101010011011111010001101100011111;
        11'd1099: TDATA = 38'b01001101001100101101100001101100011011;
        11'd1100: TDATA = 38'b01001101000101111011111001101100010101;
        11'd1101: TDATA = 38'b01001100111111001010101001101100010001;
        11'd1102: TDATA = 38'b01001100111000011001101001101100001101;
        11'd1103: TDATA = 38'b01001100110001101001000001101100001000;
        11'd1104: TDATA = 38'b01001100101010111000100001101100000100;
        11'd1105: TDATA = 38'b01001100100100001000011001101100000000;
        11'd1106: TDATA = 38'b01001100011101011000100001101011111100;
        11'd1107: TDATA = 38'b01001100010110101000111001101011111000;
        11'd1108: TDATA = 38'b01001100001111111001100001101011110011;
        11'd1109: TDATA = 38'b01001100001001001010100001101011101111;
        11'd1110: TDATA = 38'b01001100000010011011101001101011101011;
        11'd1111: TDATA = 38'b01001011111011101101001001101011100101;
        11'd1112: TDATA = 38'b01001011110100111110111001101011100001;
        11'd1113: TDATA = 38'b01001011101110010000111001101011011101;
        11'd1114: TDATA = 38'b01001011100111100011001001101011011000;
        11'd1115: TDATA = 38'b01001011100000110101110001101011010100;
        11'd1116: TDATA = 38'b01001011011010001000101001101011010000;
        11'd1117: TDATA = 38'b01001011010011011011101001101011001100;
        11'd1118: TDATA = 38'b01001011001100101111000001101011001000;
        11'd1119: TDATA = 38'b01001011000110000010110001101011000100;
        11'd1120: TDATA = 38'b01001010111111010110101001101010111111;
        11'd1121: TDATA = 38'b01001010111000101010111001101010111011;
        11'd1122: TDATA = 38'b01001010110001111111010001101010110101;
        11'd1123: TDATA = 38'b01001010101011010100000001101010110001;
        11'd1124: TDATA = 38'b01001010100100101001000001101010101101;
        11'd1125: TDATA = 38'b01001010011101111110010001101010101000;
        11'd1126: TDATA = 38'b01001010010111010011110001101010100101;
        11'd1127: TDATA = 38'b01001010010000101001101001101010100000;
        11'd1128: TDATA = 38'b01001010001001111111101001101010011100;
        11'd1129: TDATA = 38'b01001010000011010110000001101010011000;
        11'd1130: TDATA = 38'b01001001111100101100101001101010010100;
        11'd1131: TDATA = 38'b01001001110110000011100001101010010000;
        11'd1132: TDATA = 38'b01001001101111011010101001101010001100;
        11'd1133: TDATA = 38'b01001001101000110010000001101010000111;
        11'd1134: TDATA = 38'b01001001100010001001110001101010000011;
        11'd1135: TDATA = 38'b01001001011011100001101001101001111111;
        11'd1136: TDATA = 38'b01001001010100111001111001101001111001;
        11'd1137: TDATA = 38'b01001001001110010010011001101001110111;
        11'd1138: TDATA = 38'b01001001000111101011001001101001110001;
        11'd1139: TDATA = 38'b01001001000001000100001001101001101101;
        11'd1140: TDATA = 38'b01001000111010011101011001101001101001;
        11'd1141: TDATA = 38'b01001000110011110110111001101001100100;
        11'd1142: TDATA = 38'b01001000101101010000110001101001100000;
        11'd1143: TDATA = 38'b01001000100110101010110001101001011100;
        11'd1144: TDATA = 38'b01001000100000000101001001101001011000;
        11'd1145: TDATA = 38'b01001000011001011111110001101001010100;
        11'd1146: TDATA = 38'b01001000010010111010101001101001010000;
        11'd1147: TDATA = 38'b01001000001100010101110001101001001100;
        11'd1148: TDATA = 38'b01001000000101110001001001101001001000;
        11'd1149: TDATA = 38'b01000111111111001100110001101001000100;
        11'd1150: TDATA = 38'b01000111111000101000101001101000111111;
        11'd1151: TDATA = 38'b01000111110010000100111001101000111100;
        11'd1152: TDATA = 38'b01000111101011100001010001101000110111;
        11'd1153: TDATA = 38'b01000111100100111110000001101000110011;
        11'd1154: TDATA = 38'b01000111011110011011000001101000101111;
        11'd1155: TDATA = 38'b01000111010111111000001001101000101001;
        11'd1156: TDATA = 38'b01000111010001010101101001101000100101;
        11'd1157: TDATA = 38'b01000111001010110011011001101000100001;
        11'd1158: TDATA = 38'b01000111000100010001011001101000011101;
        11'd1159: TDATA = 38'b01000110111101101111101001101000011001;
        11'd1160: TDATA = 38'b01000110110111001110010001101000010101;
        11'd1161: TDATA = 38'b01000110110000101101000001101000010000;
        11'd1162: TDATA = 38'b01000110101010001100000001101000001101;
        11'd1163: TDATA = 38'b01000110100011101011011001101000001000;
        11'd1164: TDATA = 38'b01000110011101001010111001101000000100;
        11'd1165: TDATA = 38'b01000110010110101010110001101000000000;
        11'd1166: TDATA = 38'b01000110010000001010111001100111111100;
        11'd1167: TDATA = 38'b01000110001001101011001001100111111000;
        11'd1168: TDATA = 38'b01000110000011001011110001100111110100;
        11'd1169: TDATA = 38'b01000101111100101100101001100111110000;
        11'd1170: TDATA = 38'b01000101110110001101110001100111101100;
        11'd1171: TDATA = 38'b01000101101111101111001001100111101000;
        11'd1172: TDATA = 38'b01000101101001010000110001100111100100;
        11'd1173: TDATA = 38'b01000101100010110010101001100111100000;
        11'd1174: TDATA = 38'b01000101011100010100111001100111011100;
        11'd1175: TDATA = 38'b01000101010101110111010001100111010111;
        11'd1176: TDATA = 38'b01000101001111011001111001100111010100;
        11'd1177: TDATA = 38'b01000101001000111100110001100111001111;
        11'd1178: TDATA = 38'b01000101000010100000000001100111001011;
        11'd1179: TDATA = 38'b01000100111100000011011001100111001000;
        11'd1180: TDATA = 38'b01000100110101100111001001100111000011;
        11'd1181: TDATA = 38'b01000100101111001011000001100110111111;
        11'd1182: TDATA = 38'b01000100101000101111010001100110111011;
        11'd1183: TDATA = 38'b01000100100010010011110001100110110111;
        11'd1184: TDATA = 38'b01000100011011111000011001100110110011;
        11'd1185: TDATA = 38'b01000100010101011101011001100110101111;
        11'd1186: TDATA = 38'b01000100001111000010101001100110101011;
        11'd1187: TDATA = 38'b01000100001000101000000001100110100111;
        11'd1188: TDATA = 38'b01000100000010001101110001100110100011;
        11'd1189: TDATA = 38'b01000011111011110011110001100110011101;
        11'd1190: TDATA = 38'b01000011110101011010000001100110011011;
        11'd1191: TDATA = 38'b01000011101111000000100001100110010111;
        11'd1192: TDATA = 38'b01000011101000100111010001100110010001;
        11'd1193: TDATA = 38'b01000011100010001110001001100110001111;
        11'd1194: TDATA = 38'b01000011011011110101011001100110001001;
        11'd1195: TDATA = 38'b01000011010101011100111001100110000101;
        11'd1196: TDATA = 38'b01000011001111000100101001100110000011;
        11'd1197: TDATA = 38'b01000011001000101100101001100101111101;
        11'd1198: TDATA = 38'b01000011000010010100111001100101111001;
        11'd1199: TDATA = 38'b01000010111011111101011001100101110101;
        11'd1200: TDATA = 38'b01000010110101100110001001100101110001;
        11'd1201: TDATA = 38'b01000010101111001111001001100101101101;
        11'd1202: TDATA = 38'b01000010101000111000011001100101101001;
        11'd1203: TDATA = 38'b01000010100010100001111001100101100101;
        11'd1204: TDATA = 38'b01000010011100001011101001100101100001;
        11'd1205: TDATA = 38'b01000010010101110101101001100101011101;
        11'd1206: TDATA = 38'b01000010001111011111111001100101011001;
        11'd1207: TDATA = 38'b01000010001001001010011001100101010101;
        11'd1208: TDATA = 38'b01000010000010110101001001100101010001;
        11'd1209: TDATA = 38'b01000001111100100000001001100101001101;
        11'd1210: TDATA = 38'b01000001110110001011011001100101001001;
        11'd1211: TDATA = 38'b01000001101111110110111001100101000101;
        11'd1212: TDATA = 38'b01000001101001100010101001100101000001;
        11'd1213: TDATA = 38'b01000001100011001110101001100100111111;
        11'd1214: TDATA = 38'b01000001011100111010111001100100111001;
        11'd1215: TDATA = 38'b01000001010110100111011001100100110101;
        11'd1216: TDATA = 38'b01000001010000010100001001100100110011;
        11'd1217: TDATA = 38'b01000001001010000001000001100100101111;
        11'd1218: TDATA = 38'b01000001000011101110010001100100101001;
        11'd1219: TDATA = 38'b01000000111101011011110001100100100111;
        11'd1220: TDATA = 38'b01000000110111001001100001100100100011;
        11'd1221: TDATA = 38'b01000000110000110111100001100100011111;
        11'd1222: TDATA = 38'b01000000101010100101101001100100011011;
        11'd1223: TDATA = 38'b01000000100100010100001001100100010111;
        11'd1224: TDATA = 38'b01000000011110000010111001100100010011;
        11'd1225: TDATA = 38'b01000000010111110001110001100100001111;
        11'd1226: TDATA = 38'b01000000010001100001000001100100001011;
        11'd1227: TDATA = 38'b01000000001011010000011001100100000111;
        11'd1228: TDATA = 38'b01000000000101000000001001100100000100;
        11'd1229: TDATA = 38'b00111111111110110000000001100011111111;
        11'd1230: TDATA = 38'b00111111111000100000001001100011111100;
        11'd1231: TDATA = 38'b00111111110010010000101001100011111000;
        11'd1232: TDATA = 38'b00111111101100000001010001100011110100;
        11'd1233: TDATA = 38'b00111111100101110010001001100011110000;
        11'd1234: TDATA = 38'b00111111011111100011010001100011101100;
        11'd1235: TDATA = 38'b00111111011001010100101001100011101000;
        11'd1236: TDATA = 38'b00111111010011000110011001100011100100;
        11'd1237: TDATA = 38'b00111111001100111000010001100011100000;
        11'd1238: TDATA = 38'b00111111000110101010010001100011011100;
        11'd1239: TDATA = 38'b00111111000000011100101001100011011000;
        11'd1240: TDATA = 38'b00111110111010001111010001100011010100;
        11'd1241: TDATA = 38'b00111110110100000010001001100011010000;
        11'd1242: TDATA = 38'b00111110101101110101001001100011001100;
        11'd1243: TDATA = 38'b00111110100111101000100001100011001000;
        11'd1244: TDATA = 38'b00111110100001011100001001100011000100;
        11'd1245: TDATA = 38'b00111110011011001111111001100011000001;
        11'd1246: TDATA = 38'b00111110010101000011111001100010111101;
        11'd1247: TDATA = 38'b00111110001110111000010001100010111000;
        11'd1248: TDATA = 38'b00111110001000101100110001100010110101;
        11'd1249: TDATA = 38'b00111110000010100001100001100010110001;
        11'd1250: TDATA = 38'b00111101111100010110100001100010101101;
        11'd1251: TDATA = 38'b00111101110110001011110001100010101011;
        11'd1252: TDATA = 38'b00111101110000000001010001100010100111;
        11'd1253: TDATA = 38'b00111101101001110111000001100010100001;
        11'd1254: TDATA = 38'b00111101100011101100111001100010011111;
        11'd1255: TDATA = 38'b00111101011101100011001001100010011011;
        11'd1256: TDATA = 38'b00111101010111011001101001100010010111;
        11'd1257: TDATA = 38'b00111101010001010000010001100010010100;
        11'd1258: TDATA = 38'b00111101001011000111001001100010010000;
        11'd1259: TDATA = 38'b00111101000100111110011001100010001100;
        11'd1260: TDATA = 38'b00111100111110110101110001100010001000;
        11'd1261: TDATA = 38'b00111100111000101101011001100010000100;
        11'd1262: TDATA = 38'b00111100110010100101010001100010000000;
        11'd1263: TDATA = 38'b00111100101100011101010001100001111100;
        11'd1264: TDATA = 38'b00111100100110010101101001100001111000;
        11'd1265: TDATA = 38'b00111100100000001110010001100001110100;
        11'd1266: TDATA = 38'b00111100011010000111000001100001110001;
        11'd1267: TDATA = 38'b00111100010100000000001001100001101101;
        11'd1268: TDATA = 38'b00111100001101111001011001100001101001;
        11'd1269: TDATA = 38'b00111100000111110010111001100001100101;
        11'd1270: TDATA = 38'b00111100000001101100101001100001100001;
        11'd1271: TDATA = 38'b00111011111011100110101001100001011101;
        11'd1272: TDATA = 38'b00111011110101100000111001100001011011;
        11'd1273: TDATA = 38'b00111011101111011011010001100001010111;
        11'd1274: TDATA = 38'b00111011101001010110000001100001010011;
        11'd1275: TDATA = 38'b00111011100011010000111001100001010000;
        11'd1276: TDATA = 38'b00111011011101001100001001100001001100;
        11'd1277: TDATA = 38'b00111011010111000111100001100001001000;
        11'd1278: TDATA = 38'b00111011010001000011001001100001000100;
        11'd1279: TDATA = 38'b00111011001010111111000001100001000000;
        11'd1280: TDATA = 38'b00111011000100111011001001100000111100;
        11'd1281: TDATA = 38'b00111010111110110111011001100000111000;
        11'd1282: TDATA = 38'b00111010111000110100000001100000110100;
        11'd1283: TDATA = 38'b00111010110010110000110001100000110000;
        11'd1284: TDATA = 38'b00111010101100101101110001100000101101;
        11'd1285: TDATA = 38'b00111010100110101011000001100000101001;
        11'd1286: TDATA = 38'b00111010100000101000100001100000100101;
        11'd1287: TDATA = 38'b00111010011010100110010001100000100011;
        11'd1288: TDATA = 38'b00111010010100100100010001100000011111;
        11'd1289: TDATA = 38'b00111010001110100010011001100000011011;
        11'd1290: TDATA = 38'b00111010001000100000111001100000011000;
        11'd1291: TDATA = 38'b00111010000010011111100001100000010100;
        11'd1292: TDATA = 38'b00111001111100011110011001100000010000;
        11'd1293: TDATA = 38'b00111001110110011101100001100000001100;
        11'd1294: TDATA = 38'b00111001110000011100110001100000001000;
        11'd1295: TDATA = 38'b00111001101010011100011001100000000100;
        11'd1296: TDATA = 38'b00111001100100011100001001100000000001;
        11'd1297: TDATA = 38'b00111001011110011100010001011111111101;
        11'd1298: TDATA = 38'b00111001011000011100100001011111111001;
        11'd1299: TDATA = 38'b00111001010010011101000001011111110111;
        11'd1300: TDATA = 38'b00111001001100011101101001011111110011;
        11'd1301: TDATA = 38'b00111001000110011110101001011111101111;
        11'd1302: TDATA = 38'b00111001000000011111110001011111101100;
        11'd1303: TDATA = 38'b00111000111010100001010001011111101000;
        11'd1304: TDATA = 38'b00111000110100100010111001011111100100;
        11'd1305: TDATA = 38'b00111000101110100100101001011111100000;
        11'd1306: TDATA = 38'b00111000101000100110110001011111011100;
        11'd1307: TDATA = 38'b00111000100010101001001001011111011000;
        11'd1308: TDATA = 38'b00111000011100101011101001011111010101;
        11'd1309: TDATA = 38'b00111000010110101110011001011111010001;
        11'd1310: TDATA = 38'b00111000010000110001011001011111001101;
        11'd1311: TDATA = 38'b00111000001010110100101001011111001011;
        11'd1312: TDATA = 38'b00111000000100111000001001011111000111;
        11'd1313: TDATA = 38'b00110111111110111011110001011111000011;
        11'd1314: TDATA = 38'b00110111111000111111101001011111000000;
        11'd1315: TDATA = 38'b00110111110011000011110001011110111100;
        11'd1316: TDATA = 38'b00110111101101001000001001011110111000;
        11'd1317: TDATA = 38'b00110111100111001100110001011110110100;
        11'd1318: TDATA = 38'b00110111100001010001100001011110110001;
        11'd1319: TDATA = 38'b00110111011011010110101001011110101101;
        11'd1320: TDATA = 38'b00110111010101011011111001011110101001;
        11'd1321: TDATA = 38'b00110111001111100001010001011110100111;
        11'd1322: TDATA = 38'b00110111001001100111000001011110100011;
        11'd1323: TDATA = 38'b00110111000011101101000001011110011111;
        11'd1324: TDATA = 38'b00110110111101110011001001011110011100;
        11'd1325: TDATA = 38'b00110110110111111001100001011110011000;
        11'd1326: TDATA = 38'b00110110110010000000001001011110010100;
        11'd1327: TDATA = 38'b00110110101100000110111001011110010000;
        11'd1328: TDATA = 38'b00110110100110001110000001011110001101;
        11'd1329: TDATA = 38'b00110110100000010101010001011110001001;
        11'd1330: TDATA = 38'b00110110011010011100110001011110000111;
        11'd1331: TDATA = 38'b00110110010100100100100001011110000011;
        11'd1332: TDATA = 38'b00110110001110101100011001011101111111;
        11'd1333: TDATA = 38'b00110110001000110100100001011101111100;
        11'd1334: TDATA = 38'b00110110000010111100111001011101111000;
        11'd1335: TDATA = 38'b00110101111101000101100001011101110100;
        11'd1336: TDATA = 38'b00110101110111001110011001011101110000;
        11'd1337: TDATA = 38'b00110101110001010111011001011101101101;
        11'd1338: TDATA = 38'b00110101101011100000110001011101101001;
        11'd1339: TDATA = 38'b00110101100101101010010001011101100101;
        11'd1340: TDATA = 38'b00110101011111110011111001011101100011;
        11'd1341: TDATA = 38'b00110101011001111101111001011101011111;
        11'd1342: TDATA = 38'b00110101010100001000000001011101011100;
        11'd1343: TDATA = 38'b00110101001110010010011001011101011000;
        11'd1344: TDATA = 38'b00110101001000011101000001011101010100;
        11'd1345: TDATA = 38'b00110101000010100111110001011101010000;
        11'd1346: TDATA = 38'b00110100111100110010111001011101001101;
        11'd1347: TDATA = 38'b00110100110110111110001001011101001001;
        11'd1348: TDATA = 38'b00110100110001001001101001011101000111;
        11'd1349: TDATA = 38'b00110100101011010101010001011101000011;
        11'd1350: TDATA = 38'b00110100100101100001001001011101000000;
        11'd1351: TDATA = 38'b00110100011111101101011001011100111100;
        11'd1352: TDATA = 38'b00110100011001111001101001011100111000;
        11'd1353: TDATA = 38'b00110100010100000110010001011100110101;
        11'd1354: TDATA = 38'b00110100001110010011000001011100110001;
        11'd1355: TDATA = 38'b00110100001000100000000001011100101101;
        11'd1356: TDATA = 38'b00110100000010101101010001011100101011;
        11'd1357: TDATA = 38'b00110011111100111010110001011100100111;
        11'd1358: TDATA = 38'b00110011110111001000011001011100100100;
        11'd1359: TDATA = 38'b00110011110001010110010001011100100000;
        11'd1360: TDATA = 38'b00110011101011100100011001011100011100;
        11'd1361: TDATA = 38'b00110011100101110010101001011100011000;
        11'd1362: TDATA = 38'b00110011100000000001010001011100010101;
        11'd1363: TDATA = 38'b00110011011010010000000001011100010011;
        11'd1364: TDATA = 38'b00110011010100011110111001011100001111;
        11'd1365: TDATA = 38'b00110011001110101110001001011100001011;
        11'd1366: TDATA = 38'b00110011001000111101100001011100001000;
        11'd1367: TDATA = 38'b00110011000011001101001001011100000100;
        11'd1368: TDATA = 38'b00110010111101011100111001011100000000;
        11'd1369: TDATA = 38'b00110010110111101101000001011011111101;
        11'd1370: TDATA = 38'b00110010110001111101010001011011111001;
        11'd1371: TDATA = 38'b00110010101100001101110001011011110111;
        11'd1372: TDATA = 38'b00110010100110011110011001011011110011;
        11'd1373: TDATA = 38'b00110010100000101111010001011011110000;
        11'd1374: TDATA = 38'b00110010011011000000011001011011101100;
        11'd1375: TDATA = 38'b00110010010101010001110001011011101000;
        11'd1376: TDATA = 38'b00110010001111100011010001011011100101;
        11'd1377: TDATA = 38'b00110010001001110101000001011011100001;
        11'd1378: TDATA = 38'b00110010000100000111000001011011011111;
        11'd1379: TDATA = 38'b00110001111110011001010001011011011100;
        11'd1380: TDATA = 38'b00110001111000101011101001011011011000;
        11'd1381: TDATA = 38'b00110001110010111110010001011011010100;
        11'd1382: TDATA = 38'b00110001101101010001000001011011010000;
        11'd1383: TDATA = 38'b00110001100111100100001001011011001101;
        11'd1384: TDATA = 38'b00110001100001110111011001011011001001;
        11'd1385: TDATA = 38'b00110001011100001010111001011011000111;
        11'd1386: TDATA = 38'b00110001010110011110100001011011000100;
        11'd1387: TDATA = 38'b00110001010000110010011001011011000000;
        11'd1388: TDATA = 38'b00110001001011000110100001011010111100;
        11'd1389: TDATA = 38'b00110001000101011010110001011010111001;
        11'd1390: TDATA = 38'b00110000111111101111011001011010110101;
        11'd1391: TDATA = 38'b00110000111010000100000001011010110011;
        11'd1392: TDATA = 38'b00110000110100011001000001011010101111;
        11'd1393: TDATA = 38'b00110000101110101110001001011010101100;
        11'd1394: TDATA = 38'b00110000101001000011100001011010101000;
        11'd1395: TDATA = 38'b00110000100011011001001001011010100100;
        11'd1396: TDATA = 38'b00110000011101101110111001011010100001;
        11'd1397: TDATA = 38'b00110000011000000100111001011010011111;
        11'd1398: TDATA = 38'b00110000010010011011001001011010011011;
        11'd1399: TDATA = 38'b00110000001100110001100001011010011000;
        11'd1400: TDATA = 38'b00110000000111001000001001011010010100;
        11'd1401: TDATA = 38'b00110000000001011111000001011010010000;
        11'd1402: TDATA = 38'b00101111111011110110000001011010001101;
        11'd1403: TDATA = 38'b00101111110110001101011001011010001011;
        11'd1404: TDATA = 38'b00101111110000100100110001011010000111;
        11'd1405: TDATA = 38'b00101111101010111100100001011010000011;
        11'd1406: TDATA = 38'b00101111100101010100011001011010000000;
        11'd1407: TDATA = 38'b00101111011111101100100001011001111100;
        11'd1408: TDATA = 38'b00101111011010000100110001011001111001;
        11'd1409: TDATA = 38'b00101111010100011101010001011001110101;
        11'd1410: TDATA = 38'b00101111001110110110000001011001110011;
        11'd1411: TDATA = 38'b00101111001001001110111001011001110000;
        11'd1412: TDATA = 38'b00101111000011101000000001011001101100;
        11'd1413: TDATA = 38'b00101110111110000001011001011001101000;
        11'd1414: TDATA = 38'b00101110111000011010111001011001100101;
        11'd1415: TDATA = 38'b00101110110010110100101001011001100001;
        11'd1416: TDATA = 38'b00101110101101001110101001011001011111;
        11'd1417: TDATA = 38'b00101110100111101000110001011001011100;
        11'd1418: TDATA = 38'b00101110100010000011001001011001011000;
        11'd1419: TDATA = 38'b00101110011100011101110001011001010100;
        11'd1420: TDATA = 38'b00101110010110111000100001011001010001;
        11'd1421: TDATA = 38'b00101110010001010011100001011001001111;
        11'd1422: TDATA = 38'b00101110001011101110110001011001001011;
        11'd1423: TDATA = 38'b00101110000110001010001001011001001000;
        11'd1424: TDATA = 38'b00101110000000100101110001011001000100;
        11'd1425: TDATA = 38'b00101101111011000001101001011001000001;
        11'd1426: TDATA = 38'b00101101110101011101101001011000111101;
        11'd1427: TDATA = 38'b00101101101111111001110001011000111011;
        11'd1428: TDATA = 38'b00101101101010010110010001011000111000;
        11'd1429: TDATA = 38'b00101101100100110010111001011000110100;
        11'd1430: TDATA = 38'b00101101011111001111110001011000110000;
        11'd1431: TDATA = 38'b00101101011001101100110001011000101101;
        11'd1432: TDATA = 38'b00101101010100001010000001011000101011;
        11'd1433: TDATA = 38'b00101101001110100111100001011000100111;
        11'd1434: TDATA = 38'b00101101001001000101001001011000100100;
        11'd1435: TDATA = 38'b00101101000011100011000001011000100000;
        11'd1436: TDATA = 38'b00101100111110000001000001011000011101;
        11'd1437: TDATA = 38'b00101100111000011111010001011000011001;
        11'd1438: TDATA = 38'b00101100110010111101110001011000010111;
        11'd1439: TDATA = 38'b00101100101101011100011001011000010100;
        11'd1440: TDATA = 38'b00101100100111111011010001011000010000;
        11'd1441: TDATA = 38'b00101100100010011010011001011000001100;
        11'd1442: TDATA = 38'b00101100011100111001101001011000001001;
        11'd1443: TDATA = 38'b00101100010111011001001001011000000111;
        11'd1444: TDATA = 38'b00101100010001111000111001011000000011;
        11'd1445: TDATA = 38'b00101100001100011000110001011000000000;
        11'd1446: TDATA = 38'b00101100000110111000110001010111111100;
        11'd1447: TDATA = 38'b00101100000001011001001001010111111001;
        11'd1448: TDATA = 38'b00101011111011111001100001010111110111;
        11'd1449: TDATA = 38'b00101011110110011010010001010111110100;
        11'd1450: TDATA = 38'b00101011110000111011001001010111110000;
        11'd1451: TDATA = 38'b00101011101011011100010001010111101100;
        11'd1452: TDATA = 38'b00101011100101111101100001010111101001;
        11'd1453: TDATA = 38'b00101011100000011111000001010111100111;
        11'd1454: TDATA = 38'b00101011011011000000110001010111100100;
        11'd1455: TDATA = 38'b00101011010101100010101001010111100000;
        11'd1456: TDATA = 38'b00101011010000000100101001010111011100;
        11'd1457: TDATA = 38'b00101011001010100111000001010111011001;
        11'd1458: TDATA = 38'b00101011000101001001100001010111010111;
        11'd1459: TDATA = 38'b00101010111111101100001001010111010011;
        11'd1460: TDATA = 38'b00101010111010001111000001010111010000;
        11'd1461: TDATA = 38'b00101010110100110010001001010111001100;
        11'd1462: TDATA = 38'b00101010101111010101011001010111001001;
        11'd1463: TDATA = 38'b00101010101001111000111001010111000111;
        11'd1464: TDATA = 38'b00101010100100011100101001010111000100;
        11'd1465: TDATA = 38'b00101010011111000000100001010111000000;
        11'd1466: TDATA = 38'b00101010011001100100100001010110111100;
        11'd1467: TDATA = 38'b00101010010100001000111001010110111001;
        11'd1468: TDATA = 38'b00101010001110101101010001010110110111;
        11'd1469: TDATA = 38'b00101010001001010010000001010110110100;
        11'd1470: TDATA = 38'b00101010000011110110111001010110110000;
        11'd1471: TDATA = 38'b00101001111110011011111001010110101101;
        11'd1472: TDATA = 38'b00101001111001000001001001010110101011;
        11'd1473: TDATA = 38'b00101001110011100110101001010110100111;
        11'd1474: TDATA = 38'b00101001101110001100010001010110100100;
        11'd1475: TDATA = 38'b00101001101000110010001001010110100000;
        11'd1476: TDATA = 38'b00101001100011011000010001010110011101;
        11'd1477: TDATA = 38'b00101001011101111110100001010110011001;
        11'd1478: TDATA = 38'b00101001011000100100111001010110010111;
        11'd1479: TDATA = 38'b00101001010011001011100001010110010100;
        11'd1480: TDATA = 38'b00101001001101110010011001010110010000;
        11'd1481: TDATA = 38'b00101001001000011001011001010110001101;
        11'd1482: TDATA = 38'b00101001000011000000101001010110001011;
        11'd1483: TDATA = 38'b00101000111101101000000001010110001000;
        11'd1484: TDATA = 38'b00101000111000001111101001010110000100;
        11'd1485: TDATA = 38'b00101000110010110111100001010110000000;
        11'd1486: TDATA = 38'b00101000101101011111100001010101111111;
        11'd1487: TDATA = 38'b00101000101000000111101001010101111100;
        11'd1488: TDATA = 38'b00101000100010110000001001010101111000;
        11'd1489: TDATA = 38'b00101000011101011000101001010101110100;
        11'd1490: TDATA = 38'b00101000011000000001100001010101110001;
        11'd1491: TDATA = 38'b00101000010010101010011001010101101111;
        11'd1492: TDATA = 38'b00101000001101010011101001010101101100;
        11'd1493: TDATA = 38'b00101000000111111101000001010101101000;
        11'd1494: TDATA = 38'b00101000000010100110100001010101100101;
        11'd1495: TDATA = 38'b00100111111101010000010001010101100011;
        11'd1496: TDATA = 38'b00100111110111111010010001010101011111;
        11'd1497: TDATA = 38'b00100111110010100100011001010101011100;
        11'd1498: TDATA = 38'b00100111101101001110110001010101011001;
        11'd1499: TDATA = 38'b00100111100111111001010001010101010101;
        11'd1500: TDATA = 38'b00100111100010100011111001010101010011;
        11'd1501: TDATA = 38'b00100111011101001110111001010101010000;
        11'd1502: TDATA = 38'b00100111010111111010000001010101001100;
        11'd1503: TDATA = 38'b00100111010010100101010001010101001001;
        11'd1504: TDATA = 38'b00100111001101010000110001010101000111;
        11'd1505: TDATA = 38'b00100111000111111100011001010101000100;
        11'd1506: TDATA = 38'b00100111000010101000010001010101000000;
        11'd1507: TDATA = 38'b00100110111101010100011001010100111101;
        11'd1508: TDATA = 38'b00100110111000000000101001010100111011;
        11'd1509: TDATA = 38'b00100110110010101101000001010100110111;
        11'd1510: TDATA = 38'b00100110101101011001101001010100110100;
        11'd1511: TDATA = 38'b00100110101000000110100001010100110001;
        11'd1512: TDATA = 38'b00100110100010110011100001010100101101;
        11'd1513: TDATA = 38'b00100110011101100000110001010100101011;
        11'd1514: TDATA = 38'b00100110011000001110001001010100101000;
        11'd1515: TDATA = 38'b00100110010010111011101001010100100100;
        11'd1516: TDATA = 38'b00100110001101101001100001010100100001;
        11'd1517: TDATA = 38'b00100110001000010111011001010100011111;
        11'd1518: TDATA = 38'b00100110000011000101101001010100011100;
        11'd1519: TDATA = 38'b00100101111101110011111001010100011000;
        11'd1520: TDATA = 38'b00100101111000100010100001010100010101;
        11'd1521: TDATA = 38'b00100101110011010001001001010100010011;
        11'd1522: TDATA = 38'b00100101101110000000001001010100010000;
        11'd1523: TDATA = 38'b00100101101000101111001001010100001100;
        11'd1524: TDATA = 38'b00100101100011011110100001010100001001;
        11'd1525: TDATA = 38'b00100101011110001101111001010100000111;
        11'd1526: TDATA = 38'b00100101011000111101101001010100000100;
        11'd1527: TDATA = 38'b00100101010011101101100001010100000000;
        11'd1528: TDATA = 38'b00100101001110011101100001010011111101;
        11'd1529: TDATA = 38'b00100101001001001101110001010011111011;
        11'd1530: TDATA = 38'b00100101000011111110001001010011111000;
        11'd1531: TDATA = 38'b00100100111110101110110001010011110100;
        11'd1532: TDATA = 38'b00100100111001011111100001010011110001;
        11'd1533: TDATA = 38'b00100100110100010000100001010011101111;
        11'd1534: TDATA = 38'b00100100101111000001101001010011101100;
        11'd1535: TDATA = 38'b00100100101001110011000001010011101000;
        11'd1536: TDATA = 38'b00100100100100100100101001010011100101;
        11'd1537: TDATA = 38'b00100100011111010110010001010011100011;
        11'd1538: TDATA = 38'b00100100011010001000010001010011100000;
        11'd1539: TDATA = 38'b00100100010100111010010001010011011100;
        11'd1540: TDATA = 38'b00100100001111101100101001010011011001;
        11'd1541: TDATA = 38'b00100100001010011111001001010011010111;
        11'd1542: TDATA = 38'b00100100000101010001110001010011010100;
        11'd1543: TDATA = 38'b00100100000000000100101001010011010001;
        11'd1544: TDATA = 38'b00100011111010110111101001010011001101;
        11'd1545: TDATA = 38'b00100011110101101010110001010011001011;
        11'd1546: TDATA = 38'b00100011110000011110010001010011001000;
        11'd1547: TDATA = 38'b00100011101011010001110001010011000101;
        11'd1548: TDATA = 38'b00100011100110000101100001010011000011;
        11'd1549: TDATA = 38'b00100011100000111001100001010010111111;
        11'd1550: TDATA = 38'b00100011011011101101101001010010111100;
        11'd1551: TDATA = 38'b00100011010110100010000001010010111001;
        11'd1552: TDATA = 38'b00100011010001010110100001010010110111;
        11'd1553: TDATA = 38'b00100011001100001011001001010010110100;
        11'd1554: TDATA = 38'b00100011000111000000000001010010110000;
        11'd1555: TDATA = 38'b00100011000001110101001001010010101101;
        11'd1556: TDATA = 38'b00100010111100101010011001010010101011;
        11'd1557: TDATA = 38'b00100010110111011111110001010010101000;
        11'd1558: TDATA = 38'b00100010110010010101011001010010100100;
        11'd1559: TDATA = 38'b00100010101101001011001001010010100001;
        11'd1560: TDATA = 38'b00100010101000000001001001010010011111;
        11'd1561: TDATA = 38'b00100010100010110111010001010010011100;
        11'd1562: TDATA = 38'b00100010011101101101101001010010011000;
        11'd1563: TDATA = 38'b00100010011000100100001001010010010101;
        11'd1564: TDATA = 38'b00100010010011011010111001010010010100;
        11'd1565: TDATA = 38'b00100010001110010001110001010010010000;
        11'd1566: TDATA = 38'b00100010001001001000111001010010001101;
        11'd1567: TDATA = 38'b00100010000100000000001001010010001011;
        11'd1568: TDATA = 38'b00100001111110110111100001010010001000;
        11'd1569: TDATA = 38'b00100001111001101111001001010010000100;
        11'd1570: TDATA = 38'b00100001110100100110111001010010000001;
        11'd1571: TDATA = 38'b00100001101111011110111001010001111111;
        11'd1572: TDATA = 38'b00100001101010010111000001010001111100;
        11'd1573: TDATA = 38'b00100001100101001111011001010001111000;
        11'd1574: TDATA = 38'b00100001100000000111111001010001110111;
        11'd1575: TDATA = 38'b00100001011011000000101001010001110100;
        11'd1576: TDATA = 38'b00100001010101111001100001010001110000;
        11'd1577: TDATA = 38'b00100001010000110010101001010001101101;
        11'd1578: TDATA = 38'b00100001001011101011110001010001101011;
        11'd1579: TDATA = 38'b00100001000110100101010001010001101000;
        11'd1580: TDATA = 38'b00100001000001011110111001010001100100;
        11'd1581: TDATA = 38'b00100000111100011000101001010001100001;
        11'd1582: TDATA = 38'b00100000110111010010101001010001011111;
        11'd1583: TDATA = 38'b00100000110010001100110001010001011100;
        11'd1584: TDATA = 38'b00100000101101000111000001010001011001;
        11'd1585: TDATA = 38'b00100000101000000001100001010001010111;
        11'd1586: TDATA = 38'b00100000100010111100010001010001010100;
        11'd1587: TDATA = 38'b00100000011101110111001001010001010000;
        11'd1588: TDATA = 38'b00100000011000110010001001010001001101;
        11'd1589: TDATA = 38'b00100000010011101101011001010001001011;
        11'd1590: TDATA = 38'b00100000001110101000110001010001001000;
        11'd1591: TDATA = 38'b00100000001001100100011001010001000101;
        11'd1592: TDATA = 38'b00100000000100100000001001010001000011;
        11'd1593: TDATA = 38'b00011111111111011100000001010001000000;
        11'd1594: TDATA = 38'b00011111111010011000001001010000111100;
        11'd1595: TDATA = 38'b00011111110101010100011001010000111001;
        11'd1596: TDATA = 38'b00011111110000010000111001010000111000;
        11'd1597: TDATA = 38'b00011111101011001101100001010000110100;
        11'd1598: TDATA = 38'b00011111100110001010011001010000110001;
        11'd1599: TDATA = 38'b00011111100001000111011001010000101111;
        11'd1600: TDATA = 38'b00011111011100000100100001010000101100;
        11'd1601: TDATA = 38'b00011111010111000001111001010000101000;
        11'd1602: TDATA = 38'b00011111010001111111011001010000100101;
        11'd1603: TDATA = 38'b00011111001100111101001001010000100011;
        11'd1604: TDATA = 38'b00011111000111111011000001010000100000;
        11'd1605: TDATA = 38'b00011111000010111001000001010000011101;
        11'd1606: TDATA = 38'b00011110111101110111010001010000011011;
        11'd1607: TDATA = 38'b00011110111000110101101001010000011000;
        11'd1608: TDATA = 38'b00011110110011110100010001010000010100;
        11'd1609: TDATA = 38'b00011110101110110011000001010000010001;
        11'd1610: TDATA = 38'b00011110101001110001111001010000010000;
        11'd1611: TDATA = 38'b00011110100100110001000001010000001100;
        11'd1612: TDATA = 38'b00011110011111110000011001010000001001;
        11'd1613: TDATA = 38'b00011110011010101111110001010000000111;
        11'd1614: TDATA = 38'b00011110010101101111011001010000000100;
        11'd1615: TDATA = 38'b00011110010000101111010001010000000001;
        11'd1616: TDATA = 38'b00011110001011101111010001001111111111;
        11'd1617: TDATA = 38'b00011110000110101111011001001111111100;
        11'd1618: TDATA = 38'b00011110000001101111110001001111111000;
        11'd1619: TDATA = 38'b00011101111100110000010001001111110111;
        11'd1620: TDATA = 38'b00011101110111110000111001001111110100;
        11'd1621: TDATA = 38'b00011101110010110001110001001111110000;
        11'd1622: TDATA = 38'b00011101101101110010111001001111101101;
        11'd1623: TDATA = 38'b00011101101000110100000001001111101011;
        11'd1624: TDATA = 38'b00011101100011110101011001001111101000;
        11'd1625: TDATA = 38'b00011101011110110111000001001111100101;
        11'd1626: TDATA = 38'b00011101011001111000101001001111100011;
        11'd1627: TDATA = 38'b00011101010100111010101001001111100000;
        11'd1628: TDATA = 38'b00011101001111111100101001001111011100;
        11'd1629: TDATA = 38'b00011101001010111110111001001111011011;
        11'd1630: TDATA = 38'b00011101000110000001011001001111011000;
        11'd1631: TDATA = 38'b00011101000001000011111001001111010101;
        11'd1632: TDATA = 38'b00011100111100000110101001001111010011;
        11'd1633: TDATA = 38'b00011100110111001001101001001111010000;
        11'd1634: TDATA = 38'b00011100110010001100110001001111001100;
        11'd1635: TDATA = 38'b00011100101101010000000001001111001001;
        11'd1636: TDATA = 38'b00011100101000010011100001001111001000;
        11'd1637: TDATA = 38'b00011100100011010111001001001111000100;
        11'd1638: TDATA = 38'b00011100011110011010111001001111000001;
        11'd1639: TDATA = 38'b00011100011001011110111001001110111111;
        11'd1640: TDATA = 38'b00011100010100100011000001001110111100;
        11'd1641: TDATA = 38'b00011100001111100111010001001110111001;
        11'd1642: TDATA = 38'b00011100001010101011110001001110110111;
        11'd1643: TDATA = 38'b00011100000101110000011001001110110100;
        11'd1644: TDATA = 38'b00011100000000110101010001001110110001;
        11'd1645: TDATA = 38'b00011011111011111010010001001110101111;
        11'd1646: TDATA = 38'b00011011110110111111011001001110101100;
        11'd1647: TDATA = 38'b00011011110010000100110001001110101001;
        11'd1648: TDATA = 38'b00011011101101001010010001001110100111;
        11'd1649: TDATA = 38'b00011011101000001111111001001110100100;
        11'd1650: TDATA = 38'b00011011100011010101110001001110100000;
        11'd1651: TDATA = 38'b00011011011110011011110001001110011111;
        11'd1652: TDATA = 38'b00011011011001100010000001001110011100;
        11'd1653: TDATA = 38'b00011011010100101000011001001110011000;
        11'd1654: TDATA = 38'b00011011001111101110111001001110010101;
        11'd1655: TDATA = 38'b00011011001010110101100001001110010100;
        11'd1656: TDATA = 38'b00011011000101111100011001001110010000;
        11'd1657: TDATA = 38'b00011011000001000011100001001110001111;
        11'd1658: TDATA = 38'b00011010111100001010101001001110001100;
        11'd1659: TDATA = 38'b00011010110111010010000001001110001000;
        11'd1660: TDATA = 38'b00011010110010011001100001001110000101;
        11'd1661: TDATA = 38'b00011010101101100001010001001110000100;
        11'd1662: TDATA = 38'b00011010101000101001001001001110000000;
        11'd1663: TDATA = 38'b00011010100011110001001001001101111101;
        11'd1664: TDATA = 38'b00011010011110111001011001001101111011;
        11'd1665: TDATA = 38'b00011010011010000001110001001101111000;
        11'd1666: TDATA = 38'b00011010010101001010010001001101110101;
        11'd1667: TDATA = 38'b00011010010000010011000001001101110100;
        11'd1668: TDATA = 38'b00011010001011011011111001001101110000;
        11'd1669: TDATA = 38'b00011010000110100101000001001101101101;
        11'd1670: TDATA = 38'b00011010000001101110001001001101101011;
        11'd1671: TDATA = 38'b00011001111100110111100001001101101000;
        11'd1672: TDATA = 38'b00011001111000000001001001001101100101;
        11'd1673: TDATA = 38'b00011001110011001010111001001101100100;
        11'd1674: TDATA = 38'b00011001101110010100110001001101100000;
        11'd1675: TDATA = 38'b00011001101001011110110001001101011101;
        11'd1676: TDATA = 38'b00011001100100101001000001001101011011;
        11'd1677: TDATA = 38'b00011001011111110011011001001101011000;
        11'd1678: TDATA = 38'b00011001011010111101111001001101010101;
        11'd1679: TDATA = 38'b00011001010110001000101001001101010100;
        11'd1680: TDATA = 38'b00011001010001010011100001001101010000;
        11'd1681: TDATA = 38'b00011001001100011110100001001101001101;
        11'd1682: TDATA = 38'b00011001000111101001110001001101001011;
        11'd1683: TDATA = 38'b00011001000010110101001001001101001000;
        11'd1684: TDATA = 38'b00011000111110000000101001001101000101;
        11'd1685: TDATA = 38'b00011000111001001100011001001101000100;
        11'd1686: TDATA = 38'b00011000110100011000010001001101000000;
        11'd1687: TDATA = 38'b00011000101111100100010001001100111101;
        11'd1688: TDATA = 38'b00011000101010110000100001001100111011;
        11'd1689: TDATA = 38'b00011000100101111100111001001100111000;
        11'd1690: TDATA = 38'b00011000100001001001011001001100110111;
        11'd1691: TDATA = 38'b00011000011100010110001001001100110100;
        11'd1692: TDATA = 38'b00011000010111100011000001001100110000;
        11'd1693: TDATA = 38'b00011000010010110000000001001100101101;
        11'd1694: TDATA = 38'b00011000001101111101010001001100101100;
        11'd1695: TDATA = 38'b00011000001001001010100001001100101000;
        11'd1696: TDATA = 38'b00011000000100011000001001001100100111;
        11'd1697: TDATA = 38'b00010111111111100101110001001100100100;
        11'd1698: TDATA = 38'b00010111111010110011101001001100100000;
        11'd1699: TDATA = 38'b00010111110110000001101001001100011111;
        11'd1700: TDATA = 38'b00010111110001001111110001001100011100;
        11'd1701: TDATA = 38'b00010111101100011110001001001100011001;
        11'd1702: TDATA = 38'b00010111100111101100101001001100010111;
        11'd1703: TDATA = 38'b00010111100010111011010001001100010100;
        11'd1704: TDATA = 38'b00010111011110001010001001001100010001;
        11'd1705: TDATA = 38'b00010111011001011001001001001100001111;
        11'd1706: TDATA = 38'b00010111010100101000010001001100001100;
        11'd1707: TDATA = 38'b00010111001111110111100001001100001001;
        11'd1708: TDATA = 38'b00010111001011000111000001001100001000;
        11'd1709: TDATA = 38'b00010111000110010110101001001100000100;
        11'd1710: TDATA = 38'b00010111000001100110100001001100000001;
        11'd1711: TDATA = 38'b00010110111100110110011001001011111111;
        11'd1712: TDATA = 38'b00010110111000000110100001001011111100;
        11'd1713: TDATA = 38'b00010110110011010110111001001011111001;
        11'd1714: TDATA = 38'b00010110101110100111010001001011111000;
        11'd1715: TDATA = 38'b00010110101001110111111001001011110100;
        11'd1716: TDATA = 38'b00010110100101001000101001001011110011;
        11'd1717: TDATA = 38'b00010110100000011001101001001011110000;
        11'd1718: TDATA = 38'b00010110011011101010101001001011101100;
        11'd1719: TDATA = 38'b00010110010110111011111001001011101011;
        11'd1720: TDATA = 38'b00010110010010001101011001001011101000;
        11'd1721: TDATA = 38'b00010110001101011110111001001011100101;
        11'd1722: TDATA = 38'b00010110001000110000101001001011100011;
        11'd1723: TDATA = 38'b00010110000100000010100001001011100000;
        11'd1724: TDATA = 38'b00010101111111010100101001001011011101;
        11'd1725: TDATA = 38'b00010101111010100110110001001011011011;
        11'd1726: TDATA = 38'b00010101110101111001001001001011011000;
        11'd1727: TDATA = 38'b00010101110001001011101001001011010111;
        11'd1728: TDATA = 38'b00010101101100011110011001001011010100;
        11'd1729: TDATA = 38'b00010101100111110001010001001011010000;
        11'd1730: TDATA = 38'b00010101100011000100010001001011001111;
        11'd1731: TDATA = 38'b00010101011110010111011001001011001100;
        11'd1732: TDATA = 38'b00010101011001101010110001001011001001;
        11'd1733: TDATA = 38'b00010101010100111110010001001011000111;
        11'd1734: TDATA = 38'b00010101010000010001111001001011000100;
        11'd1735: TDATA = 38'b00010101001011100101101001001011000001;
        11'd1736: TDATA = 38'b00010101000110111001101001001010111111;
        11'd1737: TDATA = 38'b00010101000010001101110001001010111100;
        11'd1738: TDATA = 38'b00010100111101100010000001001010111001;
        11'd1739: TDATA = 38'b00010100111000110110100001001010111000;
        11'd1740: TDATA = 38'b00010100110100001011001001001010110101;
        11'd1741: TDATA = 38'b00010100101111011111111001001010110011;
        11'd1742: TDATA = 38'b00010100101010110100110001001010110000;
        11'd1743: TDATA = 38'b00010100100110001001111001001010101101;
        11'd1744: TDATA = 38'b00010100100001011111000001001010101011;
        11'd1745: TDATA = 38'b00010100011100110100100001001010101000;
        11'd1746: TDATA = 38'b00010100011000001010000001001010100101;
        11'd1747: TDATA = 38'b00010100010011011111110001001010100100;
        11'd1748: TDATA = 38'b00010100001110110101100001001010100000;
        11'd1749: TDATA = 38'b00010100001010001011101001001010011111;
        11'd1750: TDATA = 38'b00010100000101100001110001001010011100;
        11'd1751: TDATA = 38'b00010100000000111000001001001010011001;
        11'd1752: TDATA = 38'b00010011111100001110100001001010010111;
        11'd1753: TDATA = 38'b00010011110111100101010001001010010100;
        11'd1754: TDATA = 38'b00010011110010111100000001001010010001;
        11'd1755: TDATA = 38'b00010011101110010011000001001010010000;
        11'd1756: TDATA = 38'b00010011101001101010000001001010001100;
        11'd1757: TDATA = 38'b00010011100101000001011001001010001011;
        11'd1758: TDATA = 38'b00010011100000011000110001001010001000;
        11'd1759: TDATA = 38'b00010011011011110000011001001010000101;
        11'd1760: TDATA = 38'b00010011010111001000001001001010000011;
        11'd1761: TDATA = 38'b00010011010010100000000001001010000000;
        11'd1762: TDATA = 38'b00010011001101111000000001001001111101;
        11'd1763: TDATA = 38'b00010011001001010000010001001001111100;
        11'd1764: TDATA = 38'b00010011000100101000100001001001111000;
        11'd1765: TDATA = 38'b00010011000000000001001001001001110111;
        11'd1766: TDATA = 38'b00010010111011011001110001001001110100;
        11'd1767: TDATA = 38'b00010010110110110010101001001001110001;
        11'd1768: TDATA = 38'b00010010110010001011100001001001110000;
        11'd1769: TDATA = 38'b00010010101101100100101001001001101100;
        11'd1770: TDATA = 38'b00010010101000111110000001001001101001;
        11'd1771: TDATA = 38'b00010010100100010111011001001001101000;
        11'd1772: TDATA = 38'b00010010011111110001000001001001100100;
        11'd1773: TDATA = 38'b00010010011011001010110001001001100011;
        11'd1774: TDATA = 38'b00010010010110100100101001001001100000;
        11'd1775: TDATA = 38'b00010010010001111110110001001001011101;
        11'd1776: TDATA = 38'b00010010001101011000111001001001011100;
        11'd1777: TDATA = 38'b00010010001000110011010001001001011000;
        11'd1778: TDATA = 38'b00010010000100001101110001001001010111;
        11'd1779: TDATA = 38'b00010001111111101000100001001001010100;
        11'd1780: TDATA = 38'b00010001111011000011010001001001010001;
        11'd1781: TDATA = 38'b00010001110110011110010001001001001111;
        11'd1782: TDATA = 38'b00010001110001111001011001001001001100;
        11'd1783: TDATA = 38'b00010001101101010100101001001001001011;
        11'd1784: TDATA = 38'b00010001101000110000001001001001001000;
        11'd1785: TDATA = 38'b00010001100100001011110001001001000101;
        11'd1786: TDATA = 38'b00010001011111100111011001001001000011;
        11'd1787: TDATA = 38'b00010001011011000011011001001001000000;
        11'd1788: TDATA = 38'b00010001010110011111011001001000111101;
        11'd1789: TDATA = 38'b00010001010001111011101001001000111100;
        11'd1790: TDATA = 38'b00010001001101010111111001001000111000;
        11'd1791: TDATA = 38'b00010001001000110100011001001000110111;
        11'd1792: TDATA = 38'b00010001000100010001001001001000110100;
        11'd1793: TDATA = 38'b00010000111111101101111001001000110001;
        11'd1794: TDATA = 38'b00010000111011001010111001001000110000;
        11'd1795: TDATA = 38'b00010000110110100111111001001000101100;
        11'd1796: TDATA = 38'b00010000110010000101010001001000101011;
        11'd1797: TDATA = 38'b00010000101101100010101001001000101000;
        11'd1798: TDATA = 38'b00010000101001000000001001001000100101;
        11'd1799: TDATA = 38'b00010000100100011101111001001000100100;
        11'd1800: TDATA = 38'b00010000011111111011110001001000100000;
        11'd1801: TDATA = 38'b00010000011011011001110001001000011111;
        11'd1802: TDATA = 38'b00010000010110110111111001001000011100;
        11'd1803: TDATA = 38'b00010000010010010110010001001000011001;
        11'd1804: TDATA = 38'b00010000001101110100110001001000010111;
        11'd1805: TDATA = 38'b00010000001001010011011001001000010100;
        11'd1806: TDATA = 38'b00010000000100110010001001001000010011;
        11'd1807: TDATA = 38'b00010000000000010001000001001000010000;
        11'd1808: TDATA = 38'b00001111111011110000001001001000001101;
        11'd1809: TDATA = 38'b00001111110111001111010001001000001100;
        11'd1810: TDATA = 38'b00001111110010101110101001001000001000;
        11'd1811: TDATA = 38'b00001111101110001110001001001000000111;
        11'd1812: TDATA = 38'b00001111101001101101111001001000000100;
        11'd1813: TDATA = 38'b00001111100101001101101001001000000001;
        11'd1814: TDATA = 38'b00001111100000101101101001001000000000;
        11'd1815: TDATA = 38'b00001111011100001101110001000111111100;
        11'd1816: TDATA = 38'b00001111010111101110000001000111111011;
        11'd1817: TDATA = 38'b00001111010011001110011001000111111000;
        11'd1818: TDATA = 38'b00001111001110101111000001000111110101;
        11'd1819: TDATA = 38'b00001111001010001111101001000111110100;
        11'd1820: TDATA = 38'b00001111000101110000100001000111110000;
        11'd1821: TDATA = 38'b00001111000001010001100001000111101111;
        11'd1822: TDATA = 38'b00001110111100110010101001000111101100;
        11'd1823: TDATA = 38'b00001110111000010100000001000111101001;
        11'd1824: TDATA = 38'b00001110110011110101011001000111101000;
        11'd1825: TDATA = 38'b00001110101111010111000001000111100101;
        11'd1826: TDATA = 38'b00001110101010111000110001000111100011;
        11'd1827: TDATA = 38'b00001110100110011010101001000111100000;
        11'd1828: TDATA = 38'b00001110100001111100110001000111011101;
        11'd1829: TDATA = 38'b00001110011101011110111001000111011100;
        11'd1830: TDATA = 38'b00001110011001000001010001000111011001;
        11'd1831: TDATA = 38'b00001110010100100011110001000111010111;
        11'd1832: TDATA = 38'b00001110010000000110011001000111010100;
        11'd1833: TDATA = 38'b00001110001011101001001001000111010011;
        11'd1834: TDATA = 38'b00001110000111001100000001000111010000;
        11'd1835: TDATA = 38'b00001110000010101111001001000111001101;
        11'd1836: TDATA = 38'b00001101111110010010011001000111001100;
        11'd1837: TDATA = 38'b00001101111001110101110001000111001000;
        11'd1838: TDATA = 38'b00001101110101011001010001000111000111;
        11'd1839: TDATA = 38'b00001101110000111100111001000111000100;
        11'd1840: TDATA = 38'b00001101101100100000101001000111000001;
        11'd1841: TDATA = 38'b00001101101000000100101001000111000000;
        11'd1842: TDATA = 38'b00001101100011101000110001000110111100;
        11'd1843: TDATA = 38'b00001101011111001101000001000110111011;
        11'd1844: TDATA = 38'b00001101011010110001011001000110111000;
        11'd1845: TDATA = 38'b00001101010110010101111001000110110111;
        11'd1846: TDATA = 38'b00001101010001111010100001000110110100;
        11'd1847: TDATA = 38'b00001101001101011111011001000110110001;
        11'd1848: TDATA = 38'b00001101001001000100011001000110110000;
        11'd1849: TDATA = 38'b00001101000100101001100001000110101100;
        11'd1850: TDATA = 38'b00001101000000001110110001000110101011;
        11'd1851: TDATA = 38'b00001100111011110100001001000110101000;
        11'd1852: TDATA = 38'b00001100110111011001101001000110100101;
        11'd1853: TDATA = 38'b00001100110010111111011001000110100100;
        11'd1854: TDATA = 38'b00001100101110100101010001000110100001;
        11'd1855: TDATA = 38'b00001100101010001011001001000110100000;
        11'd1856: TDATA = 38'b00001100100101110001010001000110011100;
        11'd1857: TDATA = 38'b00001100100001010111101001000110011011;
        11'd1858: TDATA = 38'b00001100011100111110000001000110011000;
        11'd1859: TDATA = 38'b00001100011000100100100001000110010101;
        11'd1860: TDATA = 38'b00001100010100001011010001000110010100;
        11'd1861: TDATA = 38'b00001100001111110010001001000110010000;
        11'd1862: TDATA = 38'b00001100001011011001001001000110001111;
        11'd1863: TDATA = 38'b00001100000111000000010001000110001100;
        11'd1864: TDATA = 38'b00001100000010100111100001000110001011;
        11'd1865: TDATA = 38'b00001011111110001111000001000110001000;
        11'd1866: TDATA = 38'b00001011111001110110100001000110000101;
        11'd1867: TDATA = 38'b00001011110101011110010001000110000100;
        11'd1868: TDATA = 38'b00001011110001000110001001000110000001;
        11'd1869: TDATA = 38'b00001011101100101110001001000101111111;
        11'd1870: TDATA = 38'b00001011101000010110010001000101111100;
        11'd1871: TDATA = 38'b00001011100011111110100001000101111001;
        11'd1872: TDATA = 38'b00001011011111100110111001000101111000;
        11'd1873: TDATA = 38'b00001011011011001111100001000101110101;
        11'd1874: TDATA = 38'b00001011010110111000010001000101110100;
        11'd1875: TDATA = 38'b00001011010010100001000001000101110000;
        11'd1876: TDATA = 38'b00001011001110001010000001000101101111;
        11'd1877: TDATA = 38'b00001011001001110011001001000101101100;
        11'd1878: TDATA = 38'b00001011000101011100100001000101101011;
        11'd1879: TDATA = 38'b00001011000001000101111001000101101000;
        11'd1880: TDATA = 38'b00001010111100101111100001000101100101;
        11'd1881: TDATA = 38'b00001010111000011001001001000101100100;
        11'd1882: TDATA = 38'b00001010110100000011000001000101100001;
        11'd1883: TDATA = 38'b00001010101111101101000001000101011111;
        11'd1884: TDATA = 38'b00001010101011010111001001000101011100;
        11'd1885: TDATA = 38'b00001010100111000001011001000101011011;
        11'd1886: TDATA = 38'b00001010100010101011110001000101011000;
        11'd1887: TDATA = 38'b00001010011110010110011001000101010101;
        11'd1888: TDATA = 38'b00001010011010000001000001000101010100;
        11'd1889: TDATA = 38'b00001010010101101011111001000101010001;
        11'd1890: TDATA = 38'b00001010010001010110111001000101010000;
        11'd1891: TDATA = 38'b00001010001101000010000001000101001101;
        11'd1892: TDATA = 38'b00001010001000101101010001000101001011;
        11'd1893: TDATA = 38'b00001010000100011000101001000101001000;
        11'd1894: TDATA = 38'b00001010000000000100001001000101000111;
        11'd1895: TDATA = 38'b00001001111011101111111001000101000100;
        11'd1896: TDATA = 38'b00001001110111011011101001000101000001;
        11'd1897: TDATA = 38'b00001001110011000111101001000101000000;
        11'd1898: TDATA = 38'b00001001101110110011110001000100111100;
        11'd1899: TDATA = 38'b00001001101010100000000001000100111011;
        11'd1900: TDATA = 38'b00001001100110001100011001000100111000;
        11'd1901: TDATA = 38'b00001001100001111000111001000100110111;
        11'd1902: TDATA = 38'b00001001011101100101100001000100110100;
        11'd1903: TDATA = 38'b00001001011001010010010001000100110011;
        11'd1904: TDATA = 38'b00001001010100111111010001000100110000;
        11'd1905: TDATA = 38'b00001001010000101100010001000100101101;
        11'd1906: TDATA = 38'b00001001001100011001100001000100101100;
        11'd1907: TDATA = 38'b00001001001000000110111001000100101001;
        11'd1908: TDATA = 38'b00001001000011110100011001000100100111;
        11'd1909: TDATA = 38'b00001000111111100010000001000100100100;
        11'd1910: TDATA = 38'b00001000111011001111110001000100100011;
        11'd1911: TDATA = 38'b00001000110110111101101001000100100000;
        11'd1912: TDATA = 38'b00001000110010101011110001000100011101;
        11'd1913: TDATA = 38'b00001000101110011001111001000100011100;
        11'd1914: TDATA = 38'b00001000101010001000010001000100011001;
        11'd1915: TDATA = 38'b00001000100101110110101001000100011000;
        11'd1916: TDATA = 38'b00001000100001100101010001000100010101;
        11'd1917: TDATA = 38'b00001000011101010100000001000100010011;
        11'd1918: TDATA = 38'b00001000011001000010111001000100010000;
        11'd1919: TDATA = 38'b00001000010100110001111001000100001111;
        11'd1920: TDATA = 38'b00001000010000100001000001000100001100;
        11'd1921: TDATA = 38'b00001000001100010000011001000100001011;
        11'd1922: TDATA = 38'b00001000000111111111110001000100001000;
        11'd1923: TDATA = 38'b00001000000011101111010001000100000101;
        11'd1924: TDATA = 38'b00000111111111011111000001000100000100;
        11'd1925: TDATA = 38'b00000111111011001110111001000100000001;
        11'd1926: TDATA = 38'b00000111110110111110110001000011111111;
        11'd1927: TDATA = 38'b00000111110010101110111001000011111100;
        11'd1928: TDATA = 38'b00000111101110011111001001000011111011;
        11'd1929: TDATA = 38'b00000111101010001111100001000011111000;
        11'd1930: TDATA = 38'b00000111100110000000001001000011110111;
        11'd1931: TDATA = 38'b00000111100001110000110001000011110100;
        11'd1932: TDATA = 38'b00000111011101100001100001000011110001;
        11'd1933: TDATA = 38'b00000111011001010010100001000011110000;
        11'd1934: TDATA = 38'b00000111010101000011100001000011101101;
        11'd1935: TDATA = 38'b00000111010000110100110001000011101100;
        11'd1936: TDATA = 38'b00000111001100100110000001000011101001;
        11'd1937: TDATA = 38'b00000111001000010111100001000011101000;
        11'd1938: TDATA = 38'b00000111000100001001001001000011100101;
        11'd1939: TDATA = 38'b00000110111111111010111001000011100011;
        11'd1940: TDATA = 38'b00000110111011101100110001000011100000;
        11'd1941: TDATA = 38'b00000110110111011110110001000011011111;
        11'd1942: TDATA = 38'b00000110110011010000111001000011011100;
        11'd1943: TDATA = 38'b00000110101111000011010001000011011011;
        11'd1944: TDATA = 38'b00000110101010110101101001000011011000;
        11'd1945: TDATA = 38'b00000110100110101000001001000011010101;
        11'd1946: TDATA = 38'b00000110100010011010111001000011010100;
        11'd1947: TDATA = 38'b00000110011110001101101001000011010001;
        11'd1948: TDATA = 38'b00000110011010000000101001000011010000;
        11'd1949: TDATA = 38'b00000110010101110011110001000011001101;
        11'd1950: TDATA = 38'b00000110010001100111000001000011001011;
        11'd1951: TDATA = 38'b00000110001101011010011001000011001000;
        11'd1952: TDATA = 38'b00000110001001001101111001000011000111;
        11'd1953: TDATA = 38'b00000110000101000001100001000011000100;
        11'd1954: TDATA = 38'b00000110000000110101010001000011000011;
        11'd1955: TDATA = 38'b00000101111100101001001001000011000000;
        11'd1956: TDATA = 38'b00000101111000011101001001000010111111;
        11'd1957: TDATA = 38'b00000101110100010001011001000010111100;
        11'd1958: TDATA = 38'b00000101110000000101101001000010111011;
        11'd1959: TDATA = 38'b00000101101011111010000001000010111000;
        11'd1960: TDATA = 38'b00000101100111101110101001000010110101;
        11'd1961: TDATA = 38'b00000101100011100011011001000010110100;
        11'd1962: TDATA = 38'b00000101011111011000001001000010110001;
        11'd1963: TDATA = 38'b00000101011011001101001001000010110000;
        11'd1964: TDATA = 38'b00000101010111000010010001000010101101;
        11'd1965: TDATA = 38'b00000101010010110111100001000010101011;
        11'd1966: TDATA = 38'b00000101001110101100111001000010101000;
        11'd1967: TDATA = 38'b00000101001010100010011001000010100111;
        11'd1968: TDATA = 38'b00000101000110011000000001000010100100;
        11'd1969: TDATA = 38'b00000101000010001101110001000010100011;
        11'd1970: TDATA = 38'b00000100111110000011101001000010100000;
        11'd1971: TDATA = 38'b00000100111001111001101001000010011101;
        11'd1972: TDATA = 38'b00000100110101101111111001000010011100;
        11'd1973: TDATA = 38'b00000100110001100110001001000010011001;
        11'd1974: TDATA = 38'b00000100101101011100100001000010011000;
        11'd1975: TDATA = 38'b00000100101001010011001001000010010101;
        11'd1976: TDATA = 38'b00000100100101001001110001000010010100;
        11'd1977: TDATA = 38'b00000100100001000000101001000010010001;
        11'd1978: TDATA = 38'b00000100011100110111101001000010010000;
        11'd1979: TDATA = 38'b00000100011000101110101001000010001101;
        11'd1980: TDATA = 38'b00000100010100100101111001000010001100;
        11'd1981: TDATA = 38'b00000100010000011101010001000010001001;
        11'd1982: TDATA = 38'b00000100001100010100110001000010001000;
        11'd1983: TDATA = 38'b00000100001000001100011001000010000101;
        11'd1984: TDATA = 38'b00000100000100000100001001000010000100;
        11'd1985: TDATA = 38'b00000011111111111100000001000010000000;
        11'd1986: TDATA = 38'b00000011111011110100000001000001111111;
        11'd1987: TDATA = 38'b00000011110111101100001001000001111100;
        11'd1988: TDATA = 38'b00000011110011100100011001000001111011;
        11'd1989: TDATA = 38'b00000011101111011100110001000001111000;
        11'd1990: TDATA = 38'b00000011101011010101010001000001110111;
        11'd1991: TDATA = 38'b00000011100111001101111001000001110100;
        11'd1992: TDATA = 38'b00000011100011000110110001000001110011;
        11'd1993: TDATA = 38'b00000011011110111111101001000001110000;
        11'd1994: TDATA = 38'b00000011011010111000101001000001101101;
        11'd1995: TDATA = 38'b00000011010110110001111001000001101100;
        11'd1996: TDATA = 38'b00000011010010101011001001000001101001;
        11'd1997: TDATA = 38'b00000011001110100100101001000001101000;
        11'd1998: TDATA = 38'b00000011001010011110001001000001100101;
        11'd1999: TDATA = 38'b00000011000110010111111001000001100100;
        11'd2000: TDATA = 38'b00000011000010010001110001000001100001;
        11'd2001: TDATA = 38'b00000010111110001011101001000001100000;
        11'd2002: TDATA = 38'b00000010111010000101110001000001011101;
        11'd2003: TDATA = 38'b00000010110110000000000001000001011100;
        11'd2004: TDATA = 38'b00000010110001111010011001000001011000;
        11'd2005: TDATA = 38'b00000010101101110100110001000001010111;
        11'd2006: TDATA = 38'b00000010101001101111011001000001010100;
        11'd2007: TDATA = 38'b00000010100101101010001001000001010011;
        11'd2008: TDATA = 38'b00000010100001100101000001000001010000;
        11'd2009: TDATA = 38'b00000010011101100000000001000001001111;
        11'd2010: TDATA = 38'b00000010011001011011001001000001001100;
        11'd2011: TDATA = 38'b00000010010101010110011001000001001011;
        11'd2012: TDATA = 38'b00000010010001010001110001000001001000;
        11'd2013: TDATA = 38'b00000010001101001101010001000001000111;
        11'd2014: TDATA = 38'b00000010001001001000111001000001000100;
        11'd2015: TDATA = 38'b00000010000101000100101001000001000011;
        11'd2016: TDATA = 38'b00000010000001000000100001000001000000;
        11'd2017: TDATA = 38'b00000001111100111100100001000000111111;
        11'd2018: TDATA = 38'b00000001111000111000101001000000111100;
        11'd2019: TDATA = 38'b00000001110100110100111001000000111011;
        11'd2020: TDATA = 38'b00000001110000110001011001000000111000;
        11'd2021: TDATA = 38'b00000001101100101101111001000000110111;
        11'd2022: TDATA = 38'b00000001101000101010100001000000110100;
        11'd2023: TDATA = 38'b00000001100100100111010001000000110011;
        11'd2024: TDATA = 38'b00000001100000100100010001000000110000;
        11'd2025: TDATA = 38'b00000001011100100001010001000000101111;
        11'd2026: TDATA = 38'b00000001011000011110011001000000101100;
        11'd2027: TDATA = 38'b00000001010100011011110001000000101011;
        11'd2028: TDATA = 38'b00000001010000011001001001000000101000;
        11'd2029: TDATA = 38'b00000001001100010110101001000000100111;
        11'd2030: TDATA = 38'b00000001001000010100011001000000100100;
        11'd2031: TDATA = 38'b00000001000100010010001001000000100011;
        11'd2032: TDATA = 38'b00000001000000010000001001000000100000;
        11'd2033: TDATA = 38'b00000000111100001110001001000000011111;
        11'd2034: TDATA = 38'b00000000111000001100010001000000011100;
        11'd2035: TDATA = 38'b00000000110100001010101001000000011011;
        11'd2036: TDATA = 38'b00000000110000001001000001000000011000;
        11'd2037: TDATA = 38'b00000000101100000111101001000000010111;
        11'd2038: TDATA = 38'b00000000101000000110010001000000010100;
        11'd2039: TDATA = 38'b00000000100100000101001001000000010011;
        11'd2040: TDATA = 38'b00000000100000000100000001000000010000;
        11'd2041: TDATA = 38'b00000000011100000011001001000000001111;
        11'd2042: TDATA = 38'b00000000011000000010010001000000001100;
        11'd2043: TDATA = 38'b00000000010100000001101001000000001011;
        11'd2044: TDATA = 38'b00000000010000000001000001000000001000;
        11'd2045: TDATA = 38'b00000000001100000000101001000000000111;
        11'd2046: TDATA = 38'b00000000001000000000010001000000000100;
        11'd2047: TDATA = 38'b00000000000100000000001001000000000011;
        endcase
    end
    endfunction

    wire sx;
    wire [7:0] ex;
    wire [22:0] mx;
    assign sx = x[31];
    assign ex = x[30:23];
    assign mx = x[22:0];

    wire [10:0] ml;
    wire [11:0] mr;
    assign ml = x[22:12];
    assign mr = x[11:0];

    wire [37:0] tdata;
    assign tdata = TDATA(ml);

    wire [22:0] a0_inv;
    wire [14:0] a02_inv;
    assign a0_inv = tdata[37:15];
    assign a02_inv = tdata[14:0];

    wire [35:0] my_extend;
    assign my_extend = {a0_inv,13'b0} - mr * a02_inv;

    wire [22:0] my;
    assign my = my_extend[35:13];

/*
    wire [7:0] ey;
    assign ey = (253 > ex) ? 253 - ex + (mx == 23'b0): 0;
*/
    wire [8:0] eya;
    assign eya = 9'd253 + (mx == 23'b0) - ex;

    wire [7:0] ey;
    assign ey = (eya[8]) ? 0: eya[7:0];

    assign y = {sx,ey,my};

endmodule

