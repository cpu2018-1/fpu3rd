module fsqrt(
    input wire [31:0] x,
    output reg [31:0] y,
    input wire clk);

    function [39:0] TDATA (
	input [9:0] INDEX
    );
    begin
	casex(INDEX)
        10'd0: TDATA = 40'b1000011110110101011010011000110001000001;
        10'd1: TDATA = 40'b1000011110010001011010000110110011010000;
        10'd2: TDATA = 40'b1000011101110011011001110111110110111100;
        10'd3: TDATA = 40'b1000011101001111011001100101111101100010;
        10'd4: TDATA = 40'b1000011100101011011001010100000110100001;
        10'd5: TDATA = 40'b1000011100001101011001000101001111110100;
        10'd6: TDATA = 40'b1000011011101001011000110011011101001001;
        10'd7: TDATA = 40'b1000011011001011011000100100101010000100;
        10'd8: TDATA = 40'b1000011010100111011000010010111011110000;
        10'd9: TDATA = 40'b1000011010001001011000000100001100010010;
        10'd10: TDATA = 40'b1000011001100101010111110010100010010011;
        10'd11: TDATA = 40'b1000011001000111010111100011110110011101;
        10'd12: TDATA = 40'b1000011000100011010111010010010000110011;
        10'd13: TDATA = 40'b1000011000000101010111000011101000100011;
        10'd14: TDATA = 40'b1000010111100001010110110010000111001110;
        10'd15: TDATA = 40'b1000010111000011010110100011100010100101;
        10'd16: TDATA = 40'b1000010110011111010110010010000101100011;
        10'd17: TDATA = 40'b1000010110000001010110000011100100100000;
        10'd18: TDATA = 40'b1000010101100011010101110101000101000100;
        10'd19: TDATA = 40'b1000010100111111010101100011101110010011;
        10'd20: TDATA = 40'b1000010100100001010101010101010010011101;
        10'd21: TDATA = 40'b1000010100000011010101000110111000001111;
        10'd22: TDATA = 40'b1000010011011111010100110101100111101101;
        10'd23: TDATA = 40'b1000010011000001010100100111010001000100;
        10'd24: TDATA = 40'b1000010010100011010100011000111100000001;
        10'd25: TDATA = 40'b1000010010000101010100001010101000100111;
        10'd26: TDATA = 40'b1000010001100001010011111001100000010000;
        10'd27: TDATA = 40'b1000010001000011010011101011010000011001;
        10'd28: TDATA = 40'b1000010000100101010011011101000010001010;
        10'd29: TDATA = 40'b1000010000000111010011001110110101100010;
        10'd30: TDATA = 40'b1000001111100011010010111101110101010011;
        10'd31: TDATA = 40'b1000001111000101010010101111101100001110;
        10'd32: TDATA = 40'b1000001110100111010010100001100100101111;
        10'd33: TDATA = 40'b1000001110001001010010010011011110111000;
        10'd34: TDATA = 40'b1000001101101011010010000101011010100111;
        10'd35: TDATA = 40'b1000001101001101010001110111010111111100;
        10'd36: TDATA = 40'b1000001100101111010001101001010110111001;
        10'd37: TDATA = 40'b1000001100001011010001011000100100100010;
        10'd38: TDATA = 40'b1000001011101101010001001010100111000000;
        10'd39: TDATA = 40'b1000001011001111010000111100101011000100;
        10'd40: TDATA = 40'b1000001010110001010000101110110000101110;
        10'd41: TDATA = 40'b1000001010010011010000100000110111111110;
        10'd42: TDATA = 40'b1000001001110101010000010011000000110101;
        10'd43: TDATA = 40'b1000001001010111010000000101001011010001;
        10'd44: TDATA = 40'b1000001000111001001111110111010111010011;
        10'd45: TDATA = 40'b1000001000011011001111101001100100111011;
        10'd46: TDATA = 40'b1000000111111101001111011011110100001000;
        10'd47: TDATA = 40'b1000000111011111001111001110000100111011;
        10'd48: TDATA = 40'b1000000111000001001111000000010111010100;
        10'd49: TDATA = 40'b1000000110100011001110110010101011010001;
        10'd50: TDATA = 40'b1000000110000101001110100101000000110100;
        10'd51: TDATA = 40'b1000000101101101001110011010000110011001;
        10'd52: TDATA = 40'b1000000101001111001110001100011110110010;
        10'd53: TDATA = 40'b1000000100110001001101111110111000110001;
        10'd54: TDATA = 40'b1000000100010011001101110001010100010100;
        10'd55: TDATA = 40'b1000000011110101001101100011110001011100;
        10'd56: TDATA = 40'b1000000011010111001101010110010000001000;
        10'd57: TDATA = 40'b1000000010111001001101001000110000011010;
        10'd58: TDATA = 40'b1000000010100001001100111101111110100011;
        10'd59: TDATA = 40'b1000000010000011001100110000100001101001;
        10'd60: TDATA = 40'b1000000001100101001100100011000110010100;
        10'd61: TDATA = 40'b1000000001000111001100010101101100100011;
        10'd62: TDATA = 40'b1000000000101001001100001000010100010110;
        10'd63: TDATA = 40'b1000000000010001001011111101101000100001;
        10'd64: TDATA = 40'b0111111111110011001011110000010011001000;
        10'd65: TDATA = 40'b0111111111010101001011100010111111010011;
        10'd66: TDATA = 40'b0111111110111101001011011000010110111110;
        10'd67: TDATA = 40'b0111111110011111001011001011000101111101;
        10'd68: TDATA = 40'b0111111110000001001010111101110110100000;
        10'd69: TDATA = 40'b0111111101100011001010110000101000100110;
        10'd70: TDATA = 40'b0111111101001011001010100110000100111111;
        10'd71: TDATA = 40'b0111111100101101001010011000111001111001;
        10'd72: TDATA = 40'b0111111100001111001010001011110000010101;
        10'd73: TDATA = 40'b0111111011110111001010000001010000001101;
        10'd74: TDATA = 40'b0111111011011001001001110100001001011101;
        10'd75: TDATA = 40'b0111111011000001001001101001101011100100;
        10'd76: TDATA = 40'b0111111010100011001001011100100111100101;
        10'd77: TDATA = 40'b0111111010000101001001001111100101001010;
        10'd78: TDATA = 40'b0111111001101101001001000101001010101110;
        10'd79: TDATA = 40'b0111111001001111001000111000001011000100;
        10'd80: TDATA = 40'b0111111000110111001000101101110010110111;
        10'd81: TDATA = 40'b0111111000011001001000100000110101111111;
        10'd82: TDATA = 40'b0111111000000001001000010110100000000000;
        10'd83: TDATA = 40'b0111110111100011001000001001100101111001;
        10'd84: TDATA = 40'b0111110111001011000111111111010010000111;
        10'd85: TDATA = 40'b0111110110101101000111110010011010110001;
        10'd86: TDATA = 40'b0111110110010101000111101000001001001101;
        10'd87: TDATA = 40'b0111110101110111000111011011010100100111;
        10'd88: TDATA = 40'b0111110101011111000111010001000101010000;
        10'd89: TDATA = 40'b0111110101000001000111000100010011011100;
        10'd90: TDATA = 40'b0111110100101001000110111010000110010001;
        10'd91: TDATA = 40'b0111110100001011000110101101010111001101;
        10'd92: TDATA = 40'b0111110011110011000110100011001100001111;
        10'd93: TDATA = 40'b0111110011011011000110011001000010010000;
        10'd94: TDATA = 40'b0111110010111101000110001100010111001001;
        10'd95: TDATA = 40'b0111110010100101000110000010001111010111;
        10'd96: TDATA = 40'b0111110010000111000101110101100110111111;
        10'd97: TDATA = 40'b0111110001101111000101101011100001011001;
        10'd98: TDATA = 40'b0111110001010111000101100001011100110000;
        10'd99: TDATA = 40'b0111110000111001000101010100111000010101;
        10'd100: TDATA = 40'b0111110000100001000101001010110101111001;
        10'd101: TDATA = 40'b0111110000001001000101000000110100011011;
        10'd102: TDATA = 40'b0111101111101011000100110100010011111100;
        10'd103: TDATA = 40'b0111101111010011000100101010010100101001;
        10'd104: TDATA = 40'b0111101110111011000100100000010110010100;
        10'd105: TDATA = 40'b0111101110100011000100010110011000111101;
        10'd106: TDATA = 40'b0111101110000101000100001001111101100111;
        10'd107: TDATA = 40'b0111101101101101000100000000000010011011;
        10'd108: TDATA = 40'b0111101101010101000011110110001000001101;
        10'd109: TDATA = 40'b0111101100111101000011101100001110111100;
        10'd110: TDATA = 40'b0111101100011111000011011111111000101110;
        10'd111: TDATA = 40'b0111101100000111000011010110000001100111;
        10'd112: TDATA = 40'b0111101011101111000011001100001011011111;
        10'd113: TDATA = 40'b0111101011010111000011000010010110010100;
        10'd114: TDATA = 40'b0111101010111111000010111000100010000110;
        10'd115: TDATA = 40'b0111101010100001000010101100010010001011;
        10'd116: TDATA = 40'b0111101010001001000010100010100000000111;
        10'd117: TDATA = 40'b0111101001110001000010011000101111000001;
        10'd118: TDATA = 40'b0111101001011001000010001110111110111000;
        10'd119: TDATA = 40'b0111101001000001000010000101001111101100;
        10'd120: TDATA = 40'b0111101000101001000001111011100001011101;
        10'd121: TDATA = 40'b0111101000010001000001110001110100001011;
        10'd122: TDATA = 40'b0111100111110011000001100101101100111010;
        10'd123: TDATA = 40'b0111100111011011000001011100000001110010;
        10'd124: TDATA = 40'b0111100111000011000001010010010111100110;
        10'd125: TDATA = 40'b0111100110101011000001001000101110010111;
        10'd126: TDATA = 40'b0111100110010011000000111111000110000101;
        10'd127: TDATA = 40'b0111100101111011000000110101011110110000;
        10'd128: TDATA = 40'b0111100101100011000000101011111000010111;
        10'd129: TDATA = 40'b0111100101001011000000100010010010111100;
        10'd130: TDATA = 40'b0111100100110011000000011000101110011101;
        10'd131: TDATA = 40'b0111100100011011000000001111001010111010;
        10'd132: TDATA = 40'b0111100100000011000000000101101000010100;
        10'd133: TDATA = 40'b0111100011101010111111111100000110101011;
        10'd134: TDATA = 40'b0111100011010010111111110010100101111110;
        10'd135: TDATA = 40'b0111100010111010111111101001000110001101;
        10'd136: TDATA = 40'b0111100010100010111111011111100111011001;
        10'd137: TDATA = 40'b0111100010001010111111010110001001100001;
        10'd138: TDATA = 40'b0111100001110010111111001100101100100101;
        10'd139: TDATA = 40'b0111100001011010111111000011010000100110;
        10'd140: TDATA = 40'b0111100001000010111110111001110101100011;
        10'd141: TDATA = 40'b0111100000101010111110110000011011011011;
        10'd142: TDATA = 40'b0111100000010010111110100111000010010000;
        10'd143: TDATA = 40'b0111011111111010111110011101101010000001;
        10'd144: TDATA = 40'b0111011111101000111110010110101000011101;
        10'd145: TDATA = 40'b0111011111010000111110001101010001110111;
        10'd146: TDATA = 40'b0111011110111000111110000011111100001101;
        10'd147: TDATA = 40'b0111011110100000111101111010100111011111;
        10'd148: TDATA = 40'b0111011110001000111101110001010011101101;
        10'd149: TDATA = 40'b0111011101110000111101101000000000110110;
        10'd150: TDATA = 40'b0111011101011000111101011110101110111011;
        10'd151: TDATA = 40'b0111011101000000111101010101011101111100;
        10'd152: TDATA = 40'b0111011100101110111101001110100001110011;
        10'd153: TDATA = 40'b0111011100010110111101000101010010011100;
        10'd154: TDATA = 40'b0111011011111110111100111100000100000001;
        10'd155: TDATA = 40'b0111011011100110111100110010110110100001;
        10'd156: TDATA = 40'b0111011011001110111100101001101001111100;
        10'd157: TDATA = 40'b0111011010111100111100100010110001001000;
        10'd158: TDATA = 40'b0111011010100100111100011001100110001011;
        10'd159: TDATA = 40'b0111011010001100111100010000011100001010;
        10'd160: TDATA = 40'b0111011001110100111100000111010011000100;
        10'd161: TDATA = 40'b0111011001100010111100000000011100110110;
        10'd162: TDATA = 40'b0111011001001010111011110111010101011000;
        10'd163: TDATA = 40'b0111011000110010111011101110001110110101;
        10'd164: TDATA = 40'b0111011000011010111011100101001001001101;
        10'd165: TDATA = 40'b0111011000001000111011011110010101100101;
        10'd166: TDATA = 40'b0111010111110000111011010101010001100100;
        10'd167: TDATA = 40'b0111010111011000111011001100001110011110;
        10'd168: TDATA = 40'b0111010111000110111011000101011100110001;
        10'd169: TDATA = 40'b0111010110101110111010111100011011010010;
        10'd170: TDATA = 40'b0111010110010110111010110011011010101110;
        10'd171: TDATA = 40'b0111010101111110111010101010011011000101;
        10'd172: TDATA = 40'b0111010101101100111010100011101011111101;
        10'd173: TDATA = 40'b0111010101010100111010011010101101111010;
        10'd174: TDATA = 40'b0111010101000010111010010011111111111111;
        10'd175: TDATA = 40'b0111010100101010111010001011000011100011;
        10'd176: TDATA = 40'b0111010100010010111010000010001000000010;
        10'd177: TDATA = 40'b0111010100000000111001111011011100000000;
        10'd178: TDATA = 40'b0111010011101000111001110010100010000101;
        10'd179: TDATA = 40'b0111010011010000111001101001101001000100;
        10'd180: TDATA = 40'b0111010010111110111001100010111110111011;
        10'd181: TDATA = 40'b0111010010100110111001011010000111100000;
        10'd182: TDATA = 40'b0111010010010100111001010011011110100011;
        10'd183: TDATA = 40'b0111010001111100111001001010101000101111;
        10'd184: TDATA = 40'b0111010001100100111001000001110011110101;
        10'd185: TDATA = 40'b0111010001010010111000111011001100110000;
        10'd186: TDATA = 40'b0111010000111010111000110010011001011100;
        10'd187: TDATA = 40'b0111010000101000111000101011110011100011;
        10'd188: TDATA = 40'b0111010000010000111000100011000001110101;
        10'd189: TDATA = 40'b0111001111111110111000011100011101001000;
        10'd190: TDATA = 40'b0111001111100110111000010011101100111111;
        10'd191: TDATA = 40'b0111001111010100111000001101001001011111;
        10'd192: TDATA = 40'b0111001110111100111000000100011010111011;
        10'd193: TDATA = 40'b0111001110101010110111111101111000100110;
        10'd194: TDATA = 40'b0111001110010010110111110101001011101000;
        10'd195: TDATA = 40'b0111001110000000110111101110101010100000;
        10'd196: TDATA = 40'b0111001101101000110111100101111111000110;
        10'd197: TDATA = 40'b0111001101010110110111011111011111001001;
        10'd198: TDATA = 40'b0111001100111110110111010110110101010101;
        10'd199: TDATA = 40'b0111001100101100110111010000010110100100;
        10'd200: TDATA = 40'b0111001100010100110111000111101110010101;
        10'd201: TDATA = 40'b0111001100000010110111000001010000101111;
        10'd202: TDATA = 40'b0111001011110000110110111010110011101001;
        10'd203: TDATA = 40'b0111001011011000110110110010001101101010;
        10'd204: TDATA = 40'b0111001011000110110110101011110001110000;
        10'd205: TDATA = 40'b0111001010101110110110100011001101010101;
        10'd206: TDATA = 40'b0111001010011100110110011100110010100110;
        10'd207: TDATA = 40'b0111001010000100110110010100001111101111;
        10'd208: TDATA = 40'b0111001001110010110110001101110110001011;
        10'd209: TDATA = 40'b0111001001100000110110000111011101001000;
        10'd210: TDATA = 40'b0111001001001000110101111110111100100000;
        10'd211: TDATA = 40'b0111001000110110110101111000100100101000;
        10'd212: TDATA = 40'b0111001000100100110101110010001101010000;
        10'd213: TDATA = 40'b0111001000001100110101101001101110110111;
        10'd214: TDATA = 40'b0111000111111010110101100011011000101001;
        10'd215: TDATA = 40'b0111000111101000110101011101000010111100;
        10'd216: TDATA = 40'b0111000111010000110101010100100110110001;
        10'd217: TDATA = 40'b0111000110111110110101001110010010001111;
        10'd218: TDATA = 40'b0111000110101100110101000111111110001100;
        10'd219: TDATA = 40'b0111000110010100110100111111100100010000;
        10'd220: TDATA = 40'b0111000110000010110100111001010001011000;
        10'd221: TDATA = 40'b0111000101110000110100110010111111000000;
        10'd222: TDATA = 40'b0111000101011000110100101010100111010001;
        10'd223: TDATA = 40'b0111000101000110110100100100010110000100;
        10'd224: TDATA = 40'b0111000100110100110100011110000101010110;
        10'd225: TDATA = 40'b0111000100011100110100010101101111110101;
        10'd226: TDATA = 40'b0111000100001010110100001111100000010001;
        10'd227: TDATA = 40'b0111000011111000110100001001010001001110;
        10'd228: TDATA = 40'b0111000011100110110100000011000010101010;
        10'd229: TDATA = 40'b0111000011001110110011111010110000000000;
        10'd230: TDATA = 40'b0111000010111100110011110100100010100110;
        10'd231: TDATA = 40'b0111000010101010110011101110010101101100;
        10'd232: TDATA = 40'b0111000010011000110011101000001001010010;
        10'd233: TDATA = 40'b0111000010000000110011011111111001100000;
        10'd234: TDATA = 40'b0111000001101110110011011001101110001111;
        10'd235: TDATA = 40'b0111000001011100110011010011100011011110;
        10'd236: TDATA = 40'b0111000001001010110011001101011001001100;
        10'd237: TDATA = 40'b0111000000111000110011000111001111011010;
        10'd238: TDATA = 40'b0111000000100000110010111111000011001001;
        10'd239: TDATA = 40'b0111000000001110110010111000111010100001;
        10'd240: TDATA = 40'b0110111111111100110010110010110010011000;
        10'd241: TDATA = 40'b0110111111101010110010101100101010101111;
        10'd242: TDATA = 40'b0110111111011000110010100110100011100101;
        10'd243: TDATA = 40'b0110111111000110110010100000011100111011;
        10'd244: TDATA = 40'b0110111110101110110010011000010100110011;
        10'd245: TDATA = 40'b0110111110011100110010010010001111010010;
        10'd246: TDATA = 40'b0110111110001010110010001100001010010000;
        10'd247: TDATA = 40'b0110111101111000110010000110000101101110;
        10'd248: TDATA = 40'b0110111101100110110010000000000001101011;
        10'd249: TDATA = 40'b0110111101010100110001111001111110001000;
        10'd250: TDATA = 40'b0110111101000010110001110011111011000100;
        10'd251: TDATA = 40'b0110111100110000110001101101111000011111;
        10'd252: TDATA = 40'b0110111100011000110001100101110101110011;
        10'd253: TDATA = 40'b0110111100000110110001011111110100010111;
        10'd254: TDATA = 40'b0110111011110100110001011001110011011010;
        10'd255: TDATA = 40'b0110111011100010110001010011110010111101;
        10'd256: TDATA = 40'b0110111011010000110001001101110010111110;
        10'd257: TDATA = 40'b0110111010111110110001000111110011011111;
        10'd258: TDATA = 40'b0110111010101100110001000001110100011111;
        10'd259: TDATA = 40'b0110111010011010110000111011110101111110;
        10'd260: TDATA = 40'b0110111010001000110000110101110111111100;
        10'd261: TDATA = 40'b0110111001110110110000101111111010011001;
        10'd262: TDATA = 40'b0110111001100100110000101001111101010110;
        10'd263: TDATA = 40'b0110111001010010110000100100000000110001;
        10'd264: TDATA = 40'b0110111001000000110000011110000100101100;
        10'd265: TDATA = 40'b0110111000101110110000011000001001000101;
        10'd266: TDATA = 40'b0110111000011100110000010010001101111101;
        10'd267: TDATA = 40'b0110111000001010110000001100010011010101;
        10'd268: TDATA = 40'b0110110111111000110000000110011001001011;
        10'd269: TDATA = 40'b0110110111100110110000000000011111100000;
        10'd270: TDATA = 40'b0110110111010100101111111010100110010100;
        10'd271: TDATA = 40'b0110110111000010101111110100101101100111;
        10'd272: TDATA = 40'b0110110110110000101111101110110101011001;
        10'd273: TDATA = 40'b0110110110011110101111101000111101101010;
        10'd274: TDATA = 40'b0110110110001100101111100011000110011001;
        10'd275: TDATA = 40'b0110110101111010101111011101001111101000;
        10'd276: TDATA = 40'b0110110101101000101111010111011001010101;
        10'd277: TDATA = 40'b0110110101010110101111010001100011100001;
        10'd278: TDATA = 40'b0110110101000100101111001011101110001011;
        10'd279: TDATA = 40'b0110110100110010101111000101111001010101;
        10'd280: TDATA = 40'b0110110100100000101111000000000100111101;
        10'd281: TDATA = 40'b0110110100001110101110111010010001000100;
        10'd282: TDATA = 40'b0110110011111100101110110100011101101001;
        10'd283: TDATA = 40'b0110110011101010101110101110101010101101;
        10'd284: TDATA = 40'b0110110011011000101110101000111000010000;
        10'd285: TDATA = 40'b0110110011000110101110100011000110010010;
        10'd286: TDATA = 40'b0110110010110100101110011101010100110010;
        10'd287: TDATA = 40'b0110110010101000101110011001011110101101;
        10'd288: TDATA = 40'b0110110010010110101110010011101110000000;
        10'd289: TDATA = 40'b0110110010000100101110001101111101110010;
        10'd290: TDATA = 40'b0110110001110010101110001000001110000010;
        10'd291: TDATA = 40'b0110110001100000101110000010011110110000;
        10'd292: TDATA = 40'b0110110001001110101101111100101111111101;
        10'd293: TDATA = 40'b0110110000111100101101110111000001101000;
        10'd294: TDATA = 40'b0110110000101010101101110001010011110010;
        10'd295: TDATA = 40'b0110110000011110101101101101100000001010;
        10'd296: TDATA = 40'b0110110000001100101101100111110011000110;
        10'd297: TDATA = 40'b0110101111111010101101100010000110100001;
        10'd298: TDATA = 40'b0110101111101000101101011100011010011010;
        10'd299: TDATA = 40'b0110101111010110101101010110101110110010;
        10'd300: TDATA = 40'b0110101111000100101101010001000011101000;
        10'd301: TDATA = 40'b0110101110110010101101001011011000111100;
        10'd302: TDATA = 40'b0110101110100110101101000111100111011011;
        10'd303: TDATA = 40'b0110101110010100101101000001111101100010;
        10'd304: TDATA = 40'b0110101110000010101100111100010100000111;
        10'd305: TDATA = 40'b0110101101110000101100110110101011001010;
        10'd306: TDATA = 40'b0110101101011110101100110001000010101011;
        10'd307: TDATA = 40'b0110101101010010101100101101010010101000;
        10'd308: TDATA = 40'b0110101101000000101100100111101010111100;
        10'd309: TDATA = 40'b0110101100101110101100100010000011101101;
        10'd310: TDATA = 40'b0110101100011100101100011100011100111110;
        10'd311: TDATA = 40'b0110101100001010101100010110110110101100;
        10'd312: TDATA = 40'b0110101011111110101100010011001000000110;
        10'd313: TDATA = 40'b0110101011101100101100001101100010100110;
        10'd314: TDATA = 40'b0110101011011010101100000111111101100101;
        10'd315: TDATA = 40'b0110101011001000101100000010011001000001;
        10'd316: TDATA = 40'b0110101010111100101011111110101011100101;
        10'd317: TDATA = 40'b0110101010101010101011111001000111110100;
        10'd318: TDATA = 40'b0110101010011000101011110011100100100000;
        10'd319: TDATA = 40'b0110101010000110101011101110000001101011;
        10'd320: TDATA = 40'b0110101001111010101011101010010101011000;
        10'd321: TDATA = 40'b0110101001101000101011100100110011010100;
        10'd322: TDATA = 40'b0110101001010110101011011111010001101110;
        10'd323: TDATA = 40'b0110101001001010101011011011100110010001;
        10'd324: TDATA = 40'b0110101000111000101011010110000101011101;
        10'd325: TDATA = 40'b0110101000100110101011010000100101000111;
        10'd326: TDATA = 40'b0110101000010100101011001011000101001111;
        10'd327: TDATA = 40'b0110101000001000101011000111011010111010;
        10'd328: TDATA = 40'b0110100111110110101011000001111011110100;
        10'd329: TDATA = 40'b0110100111100100101010111100011101001011;
        10'd330: TDATA = 40'b0110100111011000101010111000110011101011;
        10'd331: TDATA = 40'b0110100111000110101010110011010101110101;
        10'd332: TDATA = 40'b0110100110110100101010101101111000011011;
        10'd333: TDATA = 40'b0110100110101000101010101010001111110000;
        10'd334: TDATA = 40'b0110100110010110101010100100110011001001;
        10'd335: TDATA = 40'b0110100110000100101010011111010110111111;
        10'd336: TDATA = 40'b0110100101111000101010011011101111001001;
        10'd337: TDATA = 40'b0110100101100110101010010110010011110000;
        10'd338: TDATA = 40'b0110100101010100101010010000111000110101;
        10'd339: TDATA = 40'b0110100101001000101010001101010001110100;
        10'd340: TDATA = 40'b0110100100110110101010000111110111101010;
        10'd341: TDATA = 40'b0110100100101010101010000100010001001010;
        10'd342: TDATA = 40'b0110100100011000101001111110110111110010;
        10'd343: TDATA = 40'b0110100100000110101001111001011110110111;
        10'd344: TDATA = 40'b0110100011111010101001110101111001001011;
        10'd345: TDATA = 40'b0110100011101000101001110000100001000010;
        10'd346: TDATA = 40'b0110100011010110101001101011001001010110;
        10'd347: TDATA = 40'b0110100011001010101001100111100100011110;
        10'd348: TDATA = 40'b0110100010111000101001100010001101100100;
        10'd349: TDATA = 40'b0110100010101100101001011110101001001101;
        10'd350: TDATA = 40'b0110100010011010101001011001010011000011;
        10'd351: TDATA = 40'b0110100010001000101001010011111101010111;
        10'd352: TDATA = 40'b0110100001111100101001010000011001110100;
        10'd353: TDATA = 40'b0110100001101010101001001011000100111001;
        10'd354: TDATA = 40'b0110100001011110101001000111100001110111;
        10'd355: TDATA = 40'b0110100001001100101001000010001101101101;
        10'd356: TDATA = 40'b0110100001000000101000111110101011001100;
        10'd357: TDATA = 40'b0110100000101110101000111001010111110010;
        10'd358: TDATA = 40'b0110100000011100101000110100000100110110;
        10'd359: TDATA = 40'b0110100000010000101000110000100011001001;
        10'd360: TDATA = 40'b0110011111111110101000101011010000111101;
        10'd361: TDATA = 40'b0110011111110010101000100111101111110001;
        10'd362: TDATA = 40'b0110011111100000101000100010011110010110;
        10'd363: TDATA = 40'b0110011111010100101000011110111101101010;
        10'd364: TDATA = 40'b0110011111000010101000011001101101000000;
        10'd365: TDATA = 40'b0110011110110110101000010110001100110100;
        10'd366: TDATA = 40'b0110011110100100101000010000111100111011;
        10'd367: TDATA = 40'b0110011110011000101000001101011101001111;
        10'd368: TDATA = 40'b0110011110000110101000001000001110000111;
        10'd369: TDATA = 40'b0110011101111010101000000100101110111100;
        10'd370: TDATA = 40'b0110011101101000100111111111100000100011;
        10'd371: TDATA = 40'b0110011101011100100111111100000001111001;
        10'd372: TDATA = 40'b0110011101001010100111110110110100010001;
        10'd373: TDATA = 40'b0110011100111110100111110011010110000111;
        10'd374: TDATA = 40'b0110011100101100100111101110001001001111;
        10'd375: TDATA = 40'b0110011100100000100111101010101011100101;
        10'd376: TDATA = 40'b0110011100001110100111100101011111011110;
        10'd377: TDATA = 40'b0110011100000010100111100010000010010100;
        10'd378: TDATA = 40'b0110011011110000100111011100110110111101;
        10'd379: TDATA = 40'b0110011011100100100111011001011010010100;
        10'd380: TDATA = 40'b0110011011010010100111010100001111101101;
        10'd381: TDATA = 40'b0110011011000110100111010000110011100011;
        10'd382: TDATA = 40'b0110011010110100100111001011101001101101;
        10'd383: TDATA = 40'b0110011010101000100111001000001110000100;
        10'd384: TDATA = 40'b0110011010011100100111000100110010100111;
        10'd385: TDATA = 40'b0110011010001010100110111111101001110100;
        10'd386: TDATA = 40'b0110011001111110100110111100001110110111;
        10'd387: TDATA = 40'b0110011001101100100110110111000110110101;
        10'd388: TDATA = 40'b0110011001100000100110110011101100011000;
        10'd389: TDATA = 40'b0110011001001110100110101110100101000101;
        10'd390: TDATA = 40'b0110011001000010100110101011001011001001;
        10'd391: TDATA = 40'b0110011000110110100110100111110001011001;
        10'd392: TDATA = 40'b0110011000100100100110100010101011001001;
        10'd393: TDATA = 40'b0110011000011000100110011111010001111001;
        10'd394: TDATA = 40'b0110011000000110100110011010001100011001;
        10'd395: TDATA = 40'b0110010111111010100110010110110011101001;
        10'd396: TDATA = 40'b0110010111101110100110010011011011000110;
        10'd397: TDATA = 40'b0110010111011100100110001110010110101001;
        10'd398: TDATA = 40'b0110010111010000100110001010111110100101;
        10'd399: TDATA = 40'b0110010110111110100110000101111010111000;
        10'd400: TDATA = 40'b0110010110110010100110000010100011010101;
        10'd401: TDATA = 40'b0110010110100110100101111111001011111110;
        10'd402: TDATA = 40'b0110010110010100100101111010001001010011;
        10'd403: TDATA = 40'b0110010110001000100101110110110010011100;
        10'd404: TDATA = 40'b0110010101111100100101110011011011110010;
        10'd405: TDATA = 40'b0110010101101010100101101110011010001010;
        10'd406: TDATA = 40'b0110010101011110100101101011000011111111;
        10'd407: TDATA = 40'b0110010101001100100101100110000011000111;
        10'd408: TDATA = 40'b0110010101000000100101100010101101011100;
        10'd409: TDATA = 40'b0110010100110100100101011111010111111101;
        10'd410: TDATA = 40'b0110010100100010100101011010011000000111;
        10'd411: TDATA = 40'b0110010100010110100101010111000011001000;
        10'd412: TDATA = 40'b0110010100001010100101010011101110010110;
        10'd413: TDATA = 40'b0110010011111000100101001110101111100011;
        10'd414: TDATA = 40'b0110010011101100100101001011011011010000;
        10'd415: TDATA = 40'b0110010011100000100101001000000111001010;
        10'd416: TDATA = 40'b0110010011001110100101000011001001011001;
        10'd417: TDATA = 40'b0110010011000010100100111111110101110010;
        10'd418: TDATA = 40'b0110010010110110100100111100100010011000;
        10'd419: TDATA = 40'b0110010010101010100100111001001111001011;
        10'd420: TDATA = 40'b0110010010011000100100110100010010101111;
        10'd421: TDATA = 40'b0110010010001100100100110001000000000001;
        10'd422: TDATA = 40'b0110010010000000100100101101101101100000;
        10'd423: TDATA = 40'b0110010001101110100100101000110010000101;
        10'd424: TDATA = 40'b0110010001100010100100100101100000000011;
        10'd425: TDATA = 40'b0110010001010110100100100010001110001110;
        10'd426: TDATA = 40'b0110010001001010100100011110111100100101;
        10'd427: TDATA = 40'b0110010000111000100100011010000010011111;
        10'd428: TDATA = 40'b0110010000101100100100010110110001010110;
        10'd429: TDATA = 40'b0110010000100000100100010011100000011001;
        10'd430: TDATA = 40'b0110010000001110100100001110100111010101;
        10'd431: TDATA = 40'b0110010000000010100100001011010110110111;
        10'd432: TDATA = 40'b0110001111110110100100001000000110100110;
        10'd433: TDATA = 40'b0110001111101010100100000100110110100010;
        10'd434: TDATA = 40'b0110001111011000100011111111111110110010;
        10'd435: TDATA = 40'b0110001111001100100011111100101111001100;
        10'd436: TDATA = 40'b0110001111000000100011111001011111110100;
        10'd437: TDATA = 40'b0110001110110100100011110110010000100111;
        10'd438: TDATA = 40'b0110001110100010100011110001011010001100;
        10'd439: TDATA = 40'b0110001110010110100011101110001011011110;
        10'd440: TDATA = 40'b0110001110001010100011101010111100111101;
        10'd441: TDATA = 40'b0110001101111110100011100111101110101001;
        10'd442: TDATA = 40'b0110001101110010100011100100100000100001;
        10'd443: TDATA = 40'b0110001101100000100011011111101011101100;
        10'd444: TDATA = 40'b0110001101010100100011011100011110000011;
        10'd445: TDATA = 40'b0110001101001000100011011001010000100110;
        10'd446: TDATA = 40'b0110001100111100100011010110000011010110;
        10'd447: TDATA = 40'b0110001100101010100011010001001111110101;
        10'd448: TDATA = 40'b0110001100011110100011001110000011000100;
        10'd449: TDATA = 40'b0110001100010010100011001010110110011111;
        10'd450: TDATA = 40'b0110001100000110100011000111101010000111;
        10'd451: TDATA = 40'b0110001011111010100011000100011101111011;
        10'd452: TDATA = 40'b0110001011101000100010111111101100000000;
        10'd453: TDATA = 40'b0110001011011100100010111100100000010011;
        10'd454: TDATA = 40'b0110001011010000100010111001010100110010;
        10'd455: TDATA = 40'b0110001011000100100010110110001001011110;
        10'd456: TDATA = 40'b0110001010111000100010110010111110010110;
        10'd457: TDATA = 40'b0110001010101100100010101111110011011010;
        10'd458: TDATA = 40'b0110001010011010100010101011000011011000;
        10'd459: TDATA = 40'b0110001010001110100010100111111000111011;
        10'd460: TDATA = 40'b0110001010000010100010100100101110101011;
        10'd461: TDATA = 40'b0110001001110110100010100001100100100110;
        10'd462: TDATA = 40'b0110001001101010100010011110011010101110;
        10'd463: TDATA = 40'b0110001001011110100010011011010001000011;
        10'd464: TDATA = 40'b0110001001001100100010010110100010111000;
        10'd465: TDATA = 40'b0110001001000000100010010011011001101100;
        10'd466: TDATA = 40'b0110001000110100100010010000010000101011;
        10'd467: TDATA = 40'b0110001000101000100010001101000111110111;
        10'd468: TDATA = 40'b0110001000011100100010001001111111001110;
        10'd469: TDATA = 40'b0110001000010000100010000110110110110011;
        10'd470: TDATA = 40'b0110001000000100100010000011101110100011;
        10'd471: TDATA = 40'b0110000111110010100001111111000010100011;
        10'd472: TDATA = 40'b0110000111100110100001111011111010110010;
        10'd473: TDATA = 40'b0110000111011010100001111000110011001101;
        10'd474: TDATA = 40'b0110000111001110100001110101101011110101;
        10'd475: TDATA = 40'b0110000111000010100001110010100100101000;
        10'd476: TDATA = 40'b0110000110110110100001101111011101101000;
        10'd477: TDATA = 40'b0110000110101010100001101100010110110101;
        10'd478: TDATA = 40'b0110000110011110100001101001010000001101;
        10'd479: TDATA = 40'b0110000110010010100001100110001001110010;
        10'd480: TDATA = 40'b0110000110000000100001100001100000100000;
        10'd481: TDATA = 40'b0110000101110100100001011110011010100011;
        10'd482: TDATA = 40'b0110000101101000100001011011010100110010;
        10'd483: TDATA = 40'b0110000101011100100001011000001111001101;
        10'd484: TDATA = 40'b0110000101010000100001010101001001110101;
        10'd485: TDATA = 40'b0110000101000100100001010010000100101001;
        10'd486: TDATA = 40'b0110000100111000100001001110111111101001;
        10'd487: TDATA = 40'b0110000100101100100001001011111010110101;
        10'd488: TDATA = 40'b0110000100100000100001001000110110001101;
        10'd489: TDATA = 40'b0110000100010100100001000101110001110001;
        10'd490: TDATA = 40'b0110000100001000100001000010101101100010;
        10'd491: TDATA = 40'b0110000011111100100000111111101001011111;
        10'd492: TDATA = 40'b0110000011110000100000111100100101100111;
        10'd493: TDATA = 40'b0110000011100100100000111001100001111100;
        10'd494: TDATA = 40'b0110000011010010100000110100111100110010;
        10'd495: TDATA = 40'b0110000011000110100000110001111001100101;
        10'd496: TDATA = 40'b0110000010111010100000101110110110100101;
        10'd497: TDATA = 40'b0110000010101110100000101011110011110000;
        10'd498: TDATA = 40'b0110000010100010100000101000110001000111;
        10'd499: TDATA = 40'b0110000010010110100000100101101110101011;
        10'd500: TDATA = 40'b0110000010001010100000100010101100011010;
        10'd501: TDATA = 40'b0110000001111110100000011111101010010110;
        10'd502: TDATA = 40'b0110000001110010100000011100101000011110;
        10'd503: TDATA = 40'b0110000001100110100000011001100110110010;
        10'd504: TDATA = 40'b0110000001011010100000010110100101010001;
        10'd505: TDATA = 40'b0110000001001110100000010011100011111101;
        10'd506: TDATA = 40'b0110000001000010100000010000100010110101;
        10'd507: TDATA = 40'b0110000000110110100000001101100001111001;
        10'd508: TDATA = 40'b0110000000101010100000001010100001001001;
        10'd509: TDATA = 40'b0110000000011110100000000111100000100101;
        10'd510: TDATA = 40'b0110000000010010100000000100100000001101;
        10'd511: TDATA = 40'b0110000000000110100000000001100000000001;
        10'd512: TDATA = 40'b1011111111101001111111110100000000010111;
        10'd513: TDATA = 40'b1011111110111001111111011100000011010111;
        10'd514: TDATA = 40'b1011111110001001111111000100001001010111;
        10'd515: TDATA = 40'b1011111101011001111110101100010010010110;
        10'd516: TDATA = 40'b1011111100101001111110010100011110010101;
        10'd517: TDATA = 40'b1011111011111001111101111100101101010010;
        10'd518: TDATA = 40'b1011111011001001111101100100111111001111;
        10'd519: TDATA = 40'b1011111010011111111101010000010001011000;
        10'd520: TDATA = 40'b1011111001101111111100111000101000111011;
        10'd521: TDATA = 40'b1011111000111111111100100001000011011011;
        10'd522: TDATA = 40'b1011111000001111111100001001100000111010;
        10'd523: TDATA = 40'b1011110111100101111011110100111101001001;
        10'd524: TDATA = 40'b1011110110110101111011011101100000001100;
        10'd525: TDATA = 40'b1011110110000101111011000110000110001101;
        10'd526: TDATA = 40'b1011110101010101111010101110101111001011;
        10'd527: TDATA = 40'b1011110100101011111010011010010101011101;
        10'd528: TDATA = 40'b1011110011111011111010000011000011111110;
        10'd529: TDATA = 40'b1011110011001011111001101011110101011100;
        10'd530: TDATA = 40'b1011110010100001111001010111100011001001;
        10'd531: TDATA = 40'b1011110001110001111001000000011010001001;
        10'd532: TDATA = 40'b1011110001000111111000101100001100101100;
        10'd533: TDATA = 40'b1011110000010111111000010101001001001101;
        10'd534: TDATA = 40'b1011101111101101111000000001000000100100;
        10'd535: TDATA = 40'b1011101110111101110111101010000010100110;
        10'd536: TDATA = 40'b1011101110010011110111010101111110110001;
        10'd537: TDATA = 40'b1011101101100011110110111111000110010010;
        10'd538: TDATA = 40'b1011101100111001110110101011000111010001;
        10'd539: TDATA = 40'b1011101100001001110110010100010100010010;
        10'd540: TDATA = 40'b1011101011011111110110000000011010000100;
        10'd541: TDATA = 40'b1011101010110101110101101100100010000101;
        10'd542: TDATA = 40'b1011101010000101110101010101110111000111;
        10'd543: TDATA = 40'b1011101001011011110101000010000011111011;
        10'd544: TDATA = 40'b1011101000110001110100101110010010111101;
        10'd545: TDATA = 40'b1011101000000001110100010111110000000000;
        10'd546: TDATA = 40'b1011100111010111110100000100000011110011;
        10'd547: TDATA = 40'b1011100110101101110011110000011001110100;
        10'd548: TDATA = 40'b1011100110000011110011011100110010000100;
        10'd549: TDATA = 40'b1011100101011001110011001001001100100001;
        10'd550: TDATA = 40'b1011100100101001110010110010110110101000;
        10'd551: TDATA = 40'b1011100011111111110010011111010101110101;
        10'd552: TDATA = 40'b1011100011010101110010001011110111010001;
        10'd553: TDATA = 40'b1011100010101011110001111000011010111001;
        10'd554: TDATA = 40'b1011100010000001110001100101000000110000;
        10'd555: TDATA = 40'b1011100001010111110001010001101000110011;
        10'd556: TDATA = 40'b1011100000101101110000111110010011000011;
        10'd557: TDATA = 40'b1011100000000011110000101010111111100001;
        10'd558: TDATA = 40'b1011011111011001110000010111101110001011;
        10'd559: TDATA = 40'b1011011110101111110000000100011111000010;
        10'd560: TDATA = 40'b1011011110000101101111110001010010000110;
        10'd561: TDATA = 40'b1011011101011011101111011110000111010110;
        10'd562: TDATA = 40'b1011011100110001101111001010111110110011;
        10'd563: TDATA = 40'b1011011100000111101110110111111000011100;
        10'd564: TDATA = 40'b1011011011011101101110100100110100010001;
        10'd565: TDATA = 40'b1011011010110011101110010001110010010010;
        10'd566: TDATA = 40'b1011011010001001101101111110110010011111;
        10'd567: TDATA = 40'b1011011001011111101101101011110100111000;
        10'd568: TDATA = 40'b1011011000110101101101011000111001011100;
        10'd569: TDATA = 40'b1011011000001011101101000110000000001100;
        10'd570: TDATA = 40'b1011010111100111101100110101110101011010;
        10'd571: TDATA = 40'b1011010110111101101100100011000000001101;
        10'd572: TDATA = 40'b1011010110010011101100010000001101001011;
        10'd573: TDATA = 40'b1011010101101001101011111101011100010011;
        10'd574: TDATA = 40'b1011010101000101101011101101011000101110;
        10'd575: TDATA = 40'b1011010100011011101011011010101011111000;
        10'd576: TDATA = 40'b1011010011110001101011001000000001001101;
        10'd577: TDATA = 40'b1011010011000111101010110101011000101101;
        10'd578: TDATA = 40'b1011010010100011101010100101011100010010;
        10'd579: TDATA = 40'b1011010001111001101010010010110111110010;
        10'd580: TDATA = 40'b1011010001001111101010000000010101011101;
        10'd581: TDATA = 40'b1011010000101011101001110000011110010100;
        10'd582: TDATA = 40'b1011010000000001101001011110000000000000;
        10'd583: TDATA = 40'b1011001111011101101001001110001100010010;
        10'd584: TDATA = 40'b1011001110110011101000111011110001111101;
        10'd585: TDATA = 40'b1011001110001111101000101100000001101011;
        10'd586: TDATA = 40'b1011001101100101101000011001101011010101;
        10'd587: TDATA = 40'b1011001101000001101000001001111110011110;
        10'd588: TDATA = 40'b1011001100010111100111110111101100000111;
        10'd589: TDATA = 40'b1011001011110011100111101000000010101010;
        10'd590: TDATA = 40'b1011001011001001100111010101110100010001;
        10'd591: TDATA = 40'b1011001010100101100111000110001110001110;
        10'd592: TDATA = 40'b1011001001111011100110110100000011110100;
        10'd593: TDATA = 40'b1011001001010111100110100100100001001011;
        10'd594: TDATA = 40'b1011001000101101100110010010011010101110;
        10'd595: TDATA = 40'b1011001000001001100110000010111011011110;
        10'd596: TDATA = 40'b1011000111100101100101110011011101110010;
        10'd597: TDATA = 40'b1011000110111011100101100001011101000111;
        10'd598: TDATA = 40'b1011000110010111100101010010000010110100;
        10'd599: TDATA = 40'b1011000101110011100101000010101010000100;
        10'd600: TDATA = 40'b1011000101001001100100110000101111001011;
        10'd601: TDATA = 40'b1011000100100101100100100001011001110011;
        10'd602: TDATA = 40'b1011000100000001100100010010000110000000;
        10'd603: TDATA = 40'b1011000011010111100100000000010000110110;
        10'd604: TDATA = 40'b1011000010110011100011110001000000011010;
        10'd605: TDATA = 40'b1011000010001111100011100001110001100001;
        10'd606: TDATA = 40'b1011000001101011100011010010100100001100;
        10'd607: TDATA = 40'b1011000001000111100011000011011000011010;
        10'd608: TDATA = 40'b1011000000011101100010110001101100100111;
        10'd609: TDATA = 40'b1010111111111001100010100010100100001011;
        10'd610: TDATA = 40'b1010111111010101100010010011011101010011;
        10'd611: TDATA = 40'b1010111110110001100010000100010111111101;
        10'd612: TDATA = 40'b1010111110001101100001110101010100001010;
        10'd613: TDATA = 40'b1010111101101001100001100110010001111010;
        10'd614: TDATA = 40'b1010111101000101100001010111010001001101;
        10'd615: TDATA = 40'b1010111100100001100001001000010010000010;
        10'd616: TDATA = 40'b1010111011110111100000110110110100111101;
        10'd617: TDATA = 40'b1010111011010011100000100111111001000111;
        10'd618: TDATA = 40'b1010111010101111100000011000111110110100;
        10'd619: TDATA = 40'b1010111010001011100000001010000110000011;
        10'd620: TDATA = 40'b1010111001100111011111111011001110110101;
        10'd621: TDATA = 40'b1010111001000011011111101100011001001000;
        10'd622: TDATA = 40'b1010111000011111011111011101100100111101;
        10'd623: TDATA = 40'b1010110111111011011111001110110010010101;
        10'd624: TDATA = 40'b1010110111011101011111000010011110101000;
        10'd625: TDATA = 40'b1010110110111001011110110011101110110011;
        10'd626: TDATA = 40'b1010110110010101011110100101000000100000;
        10'd627: TDATA = 40'b1010110101110001011110010110010011101110;
        10'd628: TDATA = 40'b1010110101001101011110000111101000011101;
        10'd629: TDATA = 40'b1010110100101001011101111000111110101110;
        10'd630: TDATA = 40'b1010110100000101011101101010010110100001;
        10'd631: TDATA = 40'b1010110011100001011101011011101111110101;
        10'd632: TDATA = 40'b1010110010111101011101001101001010101010;
        10'd633: TDATA = 40'b1010110010011111011101000001000010001011;
        10'd634: TDATA = 40'b1010110001111011011100110010011111110010;
        10'd635: TDATA = 40'b1010110001010111011100100011111110111010;
        10'd636: TDATA = 40'b1010110000110011011100010101011111100011;
        10'd637: TDATA = 40'b1010110000010101011100001001011011111010;
        10'd638: TDATA = 40'b1010101111110001011011111010111111010101;
        10'd639: TDATA = 40'b1010101111001101011011101100100100010000;
        10'd640: TDATA = 40'b1010101110101001011011011110001010101100;
        10'd641: TDATA = 40'b1010101110001011011011010010001011111000;
        10'd642: TDATA = 40'b1010101101100111011011000011110101000101;
        10'd643: TDATA = 40'b1010101101000011011010110101011111110010;
        10'd644: TDATA = 40'b1010101100100101011010101001100100100010;
        10'd645: TDATA = 40'b1010101100000001011010011011010010000000;
        10'd646: TDATA = 40'b1010101011011101011010001101000000111110;
        10'd647: TDATA = 40'b1010101010111111011010000001001001010000;
        10'd648: TDATA = 40'b1010101010011011011001110010111010111110;
        10'd649: TDATA = 40'b1010101001110111011001100100101110001100;
        10'd650: TDATA = 40'b1010101001011001011001011000111010000010;
        10'd651: TDATA = 40'b1010101000110101011001001010101111111111;
        10'd652: TDATA = 40'b1010101000010111011000111110111110000111;
        10'd653: TDATA = 40'b1010100111110011011000110000110110110100;
        10'd654: TDATA = 40'b1010100111010101011000100101000111001110;
        10'd655: TDATA = 40'b1010100110110001011000010111000010101010;
        10'd656: TDATA = 40'b1010100110001101011000001000111111100110;
        10'd657: TDATA = 40'b1010100101101111010111111101010011100001;
        10'd658: TDATA = 40'b1010100101001011010111101111010011001100;
        10'd659: TDATA = 40'b1010100100101101010111100011101001011000;
        10'd660: TDATA = 40'b1010100100001111010111011000000000100111;
        10'd661: TDATA = 40'b1010100011101011010111001010000100001111;
        10'd662: TDATA = 40'b1010100011001101010110111110011101101111;
        10'd663: TDATA = 40'b1010100010101001010110110000100100000110;
        10'd664: TDATA = 40'b1010100010001011010110100100111111110111;
        10'd665: TDATA = 40'b1010100001100111010110010111001000111011;
        10'd666: TDATA = 40'b1010100001001001010110001011100110111101;
        10'd667: TDATA = 40'b1010100000101011010110000000000110000000;
        10'd668: TDATA = 40'b1010100000000111010101110010010011000001;
        10'd669: TDATA = 40'b1010011111101001010101100110110100010100;
        10'd670: TDATA = 40'b1010011111001011010101011011010110101010;
        10'd671: TDATA = 40'b1010011110100111010101001101100111100111;
        10'd672: TDATA = 40'b1010011110001001010101000010001100001100;
        10'd673: TDATA = 40'b1010011101101011010100110110110001110011;
        10'd674: TDATA = 40'b1010011101000111010100101001000110101011;
        10'd675: TDATA = 40'b1010011100101001010100011101101110100010;
        10'd676: TDATA = 40'b1010011100001011010100010010010111011010;
        10'd677: TDATA = 40'b1010011011100111010100000100110000001100;
        10'd678: TDATA = 40'b1010011011001001010011111001011011010100;
        10'd679: TDATA = 40'b1010011010101011010011101110000111011101;
        10'd680: TDATA = 40'b1010011010001101010011100010110100100110;
        10'd681: TDATA = 40'b1010011001101111010011010111100010110001;
        10'd682: TDATA = 40'b1010011001001011010011001010000001111010;
        10'd683: TDATA = 40'b1010011000101101010010111110110010010100;
        10'd684: TDATA = 40'b1010011000001111010010110011100011101110;
        10'd685: TDATA = 40'b1010010111110001010010101000010110001010;
        10'd686: TDATA = 40'b1010010111010011010010011101001001100110;
        10'd687: TDATA = 40'b1010010110101111010010001111101111000100;
        10'd688: TDATA = 40'b1010010110010001010010000100100100101111;
        10'd689: TDATA = 40'b1010010101110011010001111001011011011010;
        10'd690: TDATA = 40'b1010010101010101010001101110010011000110;
        10'd691: TDATA = 40'b1010010100110111010001100011001011110011;
        10'd692: TDATA = 40'b1010010100011001010001011000000101100000;
        10'd693: TDATA = 40'b1010010011111011010001001101000000001110;
        10'd694: TDATA = 40'b1010010011011101010001000001111011111100;
        10'd695: TDATA = 40'b1010010010111111010000110110111000101010;
        10'd696: TDATA = 40'b1010010010100001010000101011110110011001;
        10'd697: TDATA = 40'b1010010010000011010000100000110101001000;
        10'd698: TDATA = 40'b1010010001100101010000010101110100111000;
        10'd699: TDATA = 40'b1010010001000111010000001010110101100111;
        10'd700: TDATA = 40'b1010010000101001001111111111110111010111;
        10'd701: TDATA = 40'b1010010000001011001111110100111010000111;
        10'd702: TDATA = 40'b1010001111101101001111101001111101110111;
        10'd703: TDATA = 40'b1010001111001111001111011111000010100111;
        10'd704: TDATA = 40'b1010001110110001001111010100001000010111;
        10'd705: TDATA = 40'b1010001110010011001111001001001111000111;
        10'd706: TDATA = 40'b1010001101110101001110111110010110110111;
        10'd707: TDATA = 40'b1010001101010111001110110011011111100111;
        10'd708: TDATA = 40'b1010001100111001001110101000101001010110;
        10'd709: TDATA = 40'b1010001100011011001110011101110100000110;
        10'd710: TDATA = 40'b1010001011111101001110010010111111110101;
        10'd711: TDATA = 40'b1010001011011111001110001000001100100011;
        10'd712: TDATA = 40'b1010001011000001001101111101011010010010;
        10'd713: TDATA = 40'b1010001010100011001101110010101000111111;
        10'd714: TDATA = 40'b1010001010001011001101101010000010010010;
        10'd715: TDATA = 40'b1010001001101101001101011111010010110010;
        10'd716: TDATA = 40'b1010001001001111001101010100100100010010;
        10'd717: TDATA = 40'b1010001000110001001101001001110110110001;
        10'd718: TDATA = 40'b1010001000010011001100111111001010001111;
        10'd719: TDATA = 40'b1010000111111011001100110110100111010101;
        10'd720: TDATA = 40'b1010000111011101001100101011111100100101;
        10'd721: TDATA = 40'b1010000110111111001100100001010010110101;
        10'd722: TDATA = 40'b1010000110100001001100010110101010000011;
        10'd723: TDATA = 40'b1010000110000011001100001100000010010001;
        10'd724: TDATA = 40'b1010000101101011001100000011100011001010;
        10'd725: TDATA = 40'b1010000101001101001011111000111101001001;
        10'd726: TDATA = 40'b1010000100101111001011101110011000000111;
        10'd727: TDATA = 40'b1010000100010001001011100011110100000101;
        10'd728: TDATA = 40'b1010000011111001001011011011010111111101;
        10'd729: TDATA = 40'b1010000011011011001011010000110101101011;
        10'd730: TDATA = 40'b1010000010111101001011000110010100011000;
        10'd731: TDATA = 40'b1010000010100101001010111101111010011101;
        10'd732: TDATA = 40'b1010000010000111001010110011011010111100;
        10'd733: TDATA = 40'b1010000001101001001010101000111100011001;
        10'd734: TDATA = 40'b1010000001010001001010100000100100101010;
        10'd735: TDATA = 40'b1010000000110011001010010110000111111000;
        10'd736: TDATA = 40'b1010000000010101001010001011101100000100;
        10'd737: TDATA = 40'b1001111111111101001010000011010110100001;
        10'd738: TDATA = 40'b1001111111011111001001111000111100011110;
        10'd739: TDATA = 40'b1001111111000001001001101110100011011010;
        10'd740: TDATA = 40'b1001111110101001001001100110010000000011;
        10'd741: TDATA = 40'b1001111110001011001001011011111000101110;
        10'd742: TDATA = 40'b1001111101110011001001010011100110110001;
        10'd743: TDATA = 40'b1001111101010101001001001001010001001101;
        10'd744: TDATA = 40'b1001111100110111001000111110111100100111;
        10'd745: TDATA = 40'b1001111100011111001000110110101100110110;
        10'd746: TDATA = 40'b1001111100000001001000101100011010000000;
        10'd747: TDATA = 40'b1001111011101001001000100100001011100111;
        10'd748: TDATA = 40'b1001111011001011001000011001111010100001;
        10'd749: TDATA = 40'b1001111010110011001000010001101101100010;
        10'd750: TDATA = 40'b1001111010010101001000000111011110001100;
        10'd751: TDATA = 40'b1001111001111101000111111111010010100110;
        10'd752: TDATA = 40'b1001111001011111000111110101000100111111;
        10'd753: TDATA = 40'b1001111001000111000111101100111010110010;
        10'd754: TDATA = 40'b1001111000101001000111100010101110111011;
        10'd755: TDATA = 40'b1001111000010001000111011010100110000111;
        10'd756: TDATA = 40'b1001110111110011000111010000011011111110;
        10'd757: TDATA = 40'b1001110111011011000111001000010100100100;
        10'd758: TDATA = 40'b1001110110111101000110111110001100001010;
        10'd759: TDATA = 40'b1001110110100101000110110110000110001000;
        10'd760: TDATA = 40'b1001110110001101000110101110000000101110;
        10'd761: TDATA = 40'b1001110101101111000110100011111010110100;
        10'd762: TDATA = 40'b1001110101010111000110011011110110110011;
        10'd763: TDATA = 40'b1001110100111001000110010001110010101000;
        10'd764: TDATA = 40'b1001110100100001000110001001101111111110;
        10'd765: TDATA = 40'b1001110100001001000110000001101101111100;
        10'd766: TDATA = 40'b1001110011101011000101110111101100010001;
        10'd767: TDATA = 40'b1001110011010011000101101111101011100111;
        10'd768: TDATA = 40'b1001110010111011000101100111101011100101;
        10'd769: TDATA = 40'b1001110010011101000101011101101100011000;
        10'd770: TDATA = 40'b1001110010000101000101010101101101101110;
        10'd771: TDATA = 40'b1001110001101101000101001101101111101011;
        10'd772: TDATA = 40'b1001110001001111000101000011110010111110;
        10'd773: TDATA = 40'b1001110000110111000100111011110110010010;
        10'd774: TDATA = 40'b1001110000011111000100110011111010001110;
        10'd775: TDATA = 40'b1001110000000001000100101010000000000000;
        10'd776: TDATA = 40'b1001101111101001000100100010000101010011;
        10'd777: TDATA = 40'b1001101111010001000100011010001011001101;
        10'd778: TDATA = 40'b1001101110110011000100010000010011011101;
        10'd779: TDATA = 40'b1001101110011011000100001000011010101111;
        10'd780: TDATA = 40'b1001101110000011000100000000100010101000;
        10'd781: TDATA = 40'b1001101101101011000011111000101011001000;
        10'd782: TDATA = 40'b1001101101001101000011101110110110100111;
        10'd783: TDATA = 40'b1001101100110101000011100111000000011110;
        10'd784: TDATA = 40'b1001101100011101000011011111001010111100;
        10'd785: TDATA = 40'b1001101100000101000011010111010110000001;
        10'd786: TDATA = 40'b1001101011101101000011001111100001101100;
        10'd787: TDATA = 40'b1001101011001111000011000101110001001001;
        10'd788: TDATA = 40'b1001101010110111000010111101111110001100;
        10'd789: TDATA = 40'b1001101010011111000010110110001011110101;
        10'd790: TDATA = 40'b1001101010000111000010101110011010000101;
        10'd791: TDATA = 40'b1001101001101111000010100110101000111100;
        10'd792: TDATA = 40'b1001101001010111000010011110111000011001;
        10'd793: TDATA = 40'b1001101000111001000010010101001100100100;
        10'd794: TDATA = 40'b1001101000100001000010001101011101011000;
        10'd795: TDATA = 40'b1001101000001001000010000101101110110011;
        10'd796: TDATA = 40'b1001100111110001000001111110000000110100;
        10'd797: TDATA = 40'b1001100111011001000001110110010011011011;
        10'd798: TDATA = 40'b1001100111000001000001101110100110101010;
        10'd799: TDATA = 40'b1001100110101001000001100110111010011110;
        10'd800: TDATA = 40'b1001100110010001000001011111001110111001;
        10'd801: TDATA = 40'b1001100101110011000001010101101001010000;
        10'd802: TDATA = 40'b1001100101011011000001001101111111000010;
        10'd803: TDATA = 40'b1001100101000011000001000110010101011001;
        10'd804: TDATA = 40'b1001100100101011000000111110101100010111;
        10'd805: TDATA = 40'b1001100100010011000000110111000011111011;
        10'd806: TDATA = 40'b1001100011111011000000101111011100000110;
        10'd807: TDATA = 40'b1001100011100011000000100111110100110110;
        10'd808: TDATA = 40'b1001100011001011000000100000001110001101;
        10'd809: TDATA = 40'b1001100010110011000000011000101000001010;
        10'd810: TDATA = 40'b1001100010011011000000010001000010101110;
        10'd811: TDATA = 40'b1001100010000011000000001001011101110111;
        10'd812: TDATA = 40'b1001100001101011000000000001111001100111;
        10'd813: TDATA = 40'b1001100001010010111111111010010101111100;
        10'd814: TDATA = 40'b1001100000111010111111110010110010111000;
        10'd815: TDATA = 40'b1001100000100010111111101011010000011010;
        10'd816: TDATA = 40'b1001100000001010111111100011101110100010;
        10'd817: TDATA = 40'b1001011111110010111111011100001101001111;
        10'd818: TDATA = 40'b1001011111011010111111010100101100100011;
        10'd819: TDATA = 40'b1001011111000010111111001101001100011101;
        10'd820: TDATA = 40'b1001011110101010111111000101101100111101;
        10'd821: TDATA = 40'b1001011110010010111110111110001110000010;
        10'd822: TDATA = 40'b1001011101111010111110110110101111101110;
        10'd823: TDATA = 40'b1001011101100010111110101111010001111111;
        10'd824: TDATA = 40'b1001011101001010111110100111110100110111;
        10'd825: TDATA = 40'b1001011100111000111110100010001111011001;
        10'd826: TDATA = 40'b1001011100100000111110011010110011010010;
        10'd827: TDATA = 40'b1001011100001000111110010011010111110001;
        10'd828: TDATA = 40'b1001011011110000111110001011111100110110;
        10'd829: TDATA = 40'b1001011011011000111110000100100010100001;
        10'd830: TDATA = 40'b1001011011000000111101111101001000110010;
        10'd831: TDATA = 40'b1001011010101000111101110101101111101000;
        10'd832: TDATA = 40'b1001011010010000111101101110010111000011;
        10'd833: TDATA = 40'b1001011001111110111101101000110101000001;
        10'd834: TDATA = 40'b1001011001100110111101100001011101011110;
        10'd835: TDATA = 40'b1001011001001110111101011010000110100010;
        10'd836: TDATA = 40'b1001011000110110111101010010110000001010;
        10'd837: TDATA = 40'b1001011000011110111101001011011010011001;
        10'd838: TDATA = 40'b1001011000000110111101000100000101001101;
        10'd839: TDATA = 40'b1001010111110100111100111110100101101100;
        10'd840: TDATA = 40'b1001010111011100111100110111010001100010;
        10'd841: TDATA = 40'b1001010111000100111100101111111101111101;
        10'd842: TDATA = 40'b1001010110101100111100101000101010111101;
        10'd843: TDATA = 40'b1001010110010100111100100001011000100011;
        10'd844: TDATA = 40'b1001010110000010111100011011111011001000;
        10'd845: TDATA = 40'b1001010101101010111100010100101001101111;
        10'd846: TDATA = 40'b1001010101010010111100001101011000111100;
        10'd847: TDATA = 40'b1001010100111010111100000110001000101101;
        10'd848: TDATA = 40'b1001010100101000111100000000101100111011;
        10'd849: TDATA = 40'b1001010100010000111011111001011101101111;
        10'd850: TDATA = 40'b1001010011111000111011110010001111000111;
        10'd851: TDATA = 40'b1001010011100000111011101011000001000101;
        10'd852: TDATA = 40'b1001010011001110111011100101100110111011;
        10'd853: TDATA = 40'b1001010010110110111011011110011001111010;
        10'd854: TDATA = 40'b1001010010011110111011010111001101011110;
        10'd855: TDATA = 40'b1001010010000110111011010000000001100111;
        10'd856: TDATA = 40'b1001010001110100111011001010101001000111;
        10'd857: TDATA = 40'b1001010001011100111011000011011110010001;
        10'd858: TDATA = 40'b1001010001000100111010111100010100000000;
        10'd859: TDATA = 40'b1001010000110010111010110110111100101100;
        10'd860: TDATA = 40'b1001010000011010111010101111110011011100;
        10'd861: TDATA = 40'b1001010000000010111010101000101010110001;
        10'd862: TDATA = 40'b1001001111110000111010100011010100101001;
        10'd863: TDATA = 40'b1001001111011000111010011100001100111111;
        10'd864: TDATA = 40'b1001001111000000111010010101000101111010;
        10'd865: TDATA = 40'b1001001110101110111010001111110000111110;
        10'd866: TDATA = 40'b1001001110010110111010001000101010111001;
        10'd867: TDATA = 40'b1001001101111110111010000001100101011010;
        10'd868: TDATA = 40'b1001001101101100111001111100010001101010;
        10'd869: TDATA = 40'b1001001101010100111001110101001101001011;
        10'd870: TDATA = 40'b1001001101000010111001101111111010001100;
        10'd871: TDATA = 40'b1001001100101010111001101000110110101101;
        10'd872: TDATA = 40'b1001001100010010111001100001110011110011;
        10'd873: TDATA = 40'b1001001100000000111001011100100010000000;
        10'd874: TDATA = 40'b1001001011101000111001010101100000000110;
        10'd875: TDATA = 40'b1001001011010110111001010000001111000011;
        10'd876: TDATA = 40'b1001001010111110111001001001001110001001;
        10'd877: TDATA = 40'b1001001010101100111001000011111101110110;
        10'd878: TDATA = 40'b1001001010010100111000111100111101111101;
        10'd879: TDATA = 40'b1001001001111100111000110101111110101001;
        10'd880: TDATA = 40'b1001001001101010111000110000101111100001;
        10'd881: TDATA = 40'b1001001001010010111000101001110001001101;
        10'd882: TDATA = 40'b1001001001000000111000100100100010110110;
        10'd883: TDATA = 40'b1001001000101000111000011101100101100001;
        10'd884: TDATA = 40'b1001001000010110111000011000010111111010;
        10'd885: TDATA = 40'b1001000111111110111000010001011011100101;
        10'd886: TDATA = 40'b1001000111101100111000001100001110101110;
        10'd887: TDATA = 40'b1001000111010100111000000101010011011001;
        10'd888: TDATA = 40'b1001000111000010111000000000000111010001;
        10'd889: TDATA = 40'b1001000110101010110111111001001100111100;
        10'd890: TDATA = 40'b1001000110011000110111110100000001100101;
        10'd891: TDATA = 40'b1001000110000000110111101101001000010000;
        10'd892: TDATA = 40'b1001000101101110110111100111111101100111;
        10'd893: TDATA = 40'b1001000101010110110111100001000101010010;
        10'd894: TDATA = 40'b1001000101000100110111011011111011011010;
        10'd895: TDATA = 40'b1001000100101100110111010101000100000100;
        10'd896: TDATA = 40'b1001000100011010110111001111111010111011;
        10'd897: TDATA = 40'b1001000100000010110111001001000100100100;
        10'd898: TDATA = 40'b1001000011110000110111000011111100001011;
        10'd899: TDATA = 40'b1001000011011110110110111110110100000111;
        10'd900: TDATA = 40'b1001000011000110110110110111111111001011;
        10'd901: TDATA = 40'b1001000010110100110110110010110111110110;
        10'd902: TDATA = 40'b1001000010011100110110101100000011111001;
        10'd903: TDATA = 40'b1001000010001010110110100110111101010011;
        10'd904: TDATA = 40'b1001000001110010110110100000001010010110;
        10'd905: TDATA = 40'b1001000001100000110110011011000100100000;
        10'd906: TDATA = 40'b1001000001001110110110010101111110111110;
        10'd907: TDATA = 40'b1001000000110110110110001111001101011011;
        10'd908: TDATA = 40'b1001000000100100110110001010001000101000;
        10'd909: TDATA = 40'b1001000000001100110110000011011000000100;
        10'd910: TDATA = 40'b1000111111111010110101111110010100000001;
        10'd911: TDATA = 40'b1000111111101000110101111001010000010001;
        10'd912: TDATA = 40'b1000111111010000110101110010100001000111;
        10'd913: TDATA = 40'b1000111110111110110101101101011110001000;
        10'd914: TDATA = 40'b1000111110101100110101101000011011011100;
        10'd915: TDATA = 40'b1000111110010100110101100001101101101100;
        10'd916: TDATA = 40'b1000111110000010110101011100101011101111;
        10'd917: TDATA = 40'b1000111101110000110101010111101010000111;
        10'd918: TDATA = 40'b1000111101011000110101010000111101110000;
        10'd919: TDATA = 40'b1000111101000110110101001011111100110111;
        10'd920: TDATA = 40'b1000111100110100110101000110111100010010;
        10'd921: TDATA = 40'b1000111100011100110101000000010001010101;
        10'd922: TDATA = 40'b1000111100001010110100111011010001011110;
        10'd923: TDATA = 40'b1000111011111000110100110110010001111100;
        10'd924: TDATA = 40'b1000111011100000110100101111101000011001;
        10'd925: TDATA = 40'b1000111011001110110100101010101001100110;
        10'd926: TDATA = 40'b1000111010111100110100100101101011000110;
        10'd927: TDATA = 40'b1000111010101010110100100000101100111011;
        10'd928: TDATA = 40'b1000111010010010110100011010000101001100;
        10'd929: TDATA = 40'b1000111010000000110100010101000111110000;
        10'd930: TDATA = 40'b1000111001101110110100010000001010100111;
        10'd931: TDATA = 40'b1000111001010110110100001001100100010001;
        10'd932: TDATA = 40'b1000111001000100110100000100100111110111;
        10'd933: TDATA = 40'b1000111000110010110011111111101011110010;
        10'd934: TDATA = 40'b1000111000100000110011111010110000000000;
        10'd935: TDATA = 40'b1000111000001000110011110100001011011101;
        10'd936: TDATA = 40'b1000110111110110110011101111010000011010;
        10'd937: TDATA = 40'b1000110111100100110011101010010101101100;
        10'd938: TDATA = 40'b1000110111010010110011100101011011010001;
        10'd939: TDATA = 40'b1000110111000000110011100000100001001010;
        10'd940: TDATA = 40'b1000110110101000110011011001111110110100;
        10'd941: TDATA = 40'b1000110110010110110011010101000101011100;
        10'd942: TDATA = 40'b1000110110000100110011010000001100010111;
        10'd943: TDATA = 40'b1000110101110010110011001011010011100111;
        10'd944: TDATA = 40'b1000110101011010110011000100110011000101;
        10'd945: TDATA = 40'b1000110101001000110010111111111011000010;
        10'd946: TDATA = 40'b1000110100110110110010111011000011010100;
        10'd947: TDATA = 40'b1000110100100100110010110110001011111001;
        10'd948: TDATA = 40'b1000110100010010110010110001010100110010;
        10'd949: TDATA = 40'b1000110100000000110010101100011110000000;
        10'd950: TDATA = 40'b1000110011101000110010100110000000000101;
        10'd951: TDATA = 40'b1000110011010110110010100001001010000000;
        10'd952: TDATA = 40'b1000110011000100110010011100010100010000;
        10'd953: TDATA = 40'b1000110010110010110010010111011110110011;
        10'd954: TDATA = 40'b1000110010100000110010010010101001101001;
        10'd955: TDATA = 40'b1000110010001110110010001101110100110100;
        10'd956: TDATA = 40'b1000110001111100110010001001000000010010;
        10'd957: TDATA = 40'b1000110001100100110010000010100101011001;
        10'd958: TDATA = 40'b1000110001010010110001111101110001100101;
        10'd959: TDATA = 40'b1000110001000000110001111000111110000110;
        10'd960: TDATA = 40'b1000110000101110110001110100001010111001;
        10'd961: TDATA = 40'b1000110000011100110001101111011000000001;
        10'd962: TDATA = 40'b1000110000001010110001101010100101011100;
        10'd963: TDATA = 40'b1000101111111000110001100101110011001011;
        10'd964: TDATA = 40'b1000101111100110110001100001000001001110;
        10'd965: TDATA = 40'b1000101111010100110001011100001111100100;
        10'd966: TDATA = 40'b1000101110111100110001010101111000100000;
        10'd967: TDATA = 40'b1000101110101010110001010001000111100100;
        10'd968: TDATA = 40'b1000101110011000110001001100010110111100;
        10'd969: TDATA = 40'b1000101110000110110001000111100110100111;
        10'd970: TDATA = 40'b1000101101110100110001000010110110100110;
        10'd971: TDATA = 40'b1000101101100010110000111110000110111001;
        10'd972: TDATA = 40'b1000101101010000110000111001010111011111;
        10'd973: TDATA = 40'b1000101100111110110000110100101000011001;
        10'd974: TDATA = 40'b1000101100101100110000101111111001100110;
        10'd975: TDATA = 40'b1000101100011010110000101011001011000111;
        10'd976: TDATA = 40'b1000101100001000110000100110011100111100;
        10'd977: TDATA = 40'b1000101011110110110000100001101111000100;
        10'd978: TDATA = 40'b1000101011100100110000011101000001100000;
        10'd979: TDATA = 40'b1000101011010010110000011000010100001111;
        10'd980: TDATA = 40'b1000101011000000110000010011100111010010;
        10'd981: TDATA = 40'b1000101010101110110000001110111010101000;
        10'd982: TDATA = 40'b1000101010011100110000001010001110010001;
        10'd983: TDATA = 40'b1000101010001010110000000101100010001111;
        10'd984: TDATA = 40'b1000101001111000110000000000110110011111;
        10'd985: TDATA = 40'b1000101001100110101111111100001011000011;
        10'd986: TDATA = 40'b1000101001010100101111110111011111111011;
        10'd987: TDATA = 40'b1000101001000010101111110010110101000110;
        10'd988: TDATA = 40'b1000101000110000101111101110001010100101;
        10'd989: TDATA = 40'b1000101000011110101111101001100000010110;
        10'd990: TDATA = 40'b1000101000001100101111100100110110011100;
        10'd991: TDATA = 40'b1000100111111010101111100000001100110101;
        10'd992: TDATA = 40'b1000100111101000101111011011100011100001;
        10'd993: TDATA = 40'b1000100111010110101111010110111010100000;
        10'd994: TDATA = 40'b1000100111000100101111010010010001110011;
        10'd995: TDATA = 40'b1000100110110010101111001101101001011010;
        10'd996: TDATA = 40'b1000100110100000101111001001000001010011;
        10'd997: TDATA = 40'b1000100110001110101111000100011001100000;
        10'd998: TDATA = 40'b1000100101111100101110111111110010000001;
        10'd999: TDATA = 40'b1000100101101010101110111011001010110100;
        10'd1000: TDATA = 40'b1000100101011000101110110110100011111011;
        10'd1001: TDATA = 40'b1000100101000110101110110001111101010110;
        10'd1002: TDATA = 40'b1000100100110100101110101101010111000011;
        10'd1003: TDATA = 40'b1000100100100010101110101000110001000100;
        10'd1004: TDATA = 40'b1000100100010110101110100101101101010000;
        10'd1005: TDATA = 40'b1000100100000100101110100001000111110001;
        10'd1006: TDATA = 40'b1000100011110010101110011100100010100101;
        10'd1007: TDATA = 40'b1000100011100000101110010111111101101101;
        10'd1008: TDATA = 40'b1000100011001110101110010011011001001000;
        10'd1009: TDATA = 40'b1000100010111100101110001110110100110110;
        10'd1010: TDATA = 40'b1000100010101010101110001010010000110111;
        10'd1011: TDATA = 40'b1000100010011000101110000101101101001100;
        10'd1012: TDATA = 40'b1000100010000110101110000001001001110011;
        10'd1013: TDATA = 40'b1000100001111010101101111110000111101110;
        10'd1014: TDATA = 40'b1000100001101000101101111001100100110110;
        10'd1015: TDATA = 40'b1000100001010110101101110101000010010000;
        10'd1016: TDATA = 40'b1000100001000100101101110000011111111111;
        10'd1017: TDATA = 40'b1000100000110010101101101011111110000000;
        10'd1018: TDATA = 40'b1000100000100000101101100111011100010100;
        10'd1019: TDATA = 40'b1000100000001110101101100010111010111100;
        10'd1020: TDATA = 40'b1000100000000010101101011111111010001011;
        10'd1021: TDATA = 40'b1000011111110000101101011011011001010011;
        10'd1022: TDATA = 40'b1000011111011110101101010110111000101101;
        10'd1023: TDATA = 40'b1000011111001100101101010010011000011011;
	endcase
    end
    endfunction

    reg [7:0] ey_reg1,ey_reg2,ey_reg3;
    reg [14:0] thalf_x0_reg1,thalf_x0_reg2;
    reg [22:0] mr_reg,mx_reg1,mx_reg2,mx_reg3;
    reg [23:0] half_ax03_reg;
    reg [24:0] half_x03_reg;

    // stage1
    wire odd_flag;
    wire [7:0] ex;
    wire [22:0] mx;
    wire [11:0] index;
    assign odd_flag = x[23];
    assign ex = x[30:23];
    assign mx = x[22:0];
    assign index = x[23:14];

    wire [39:0] tdata;
    assign tdata = TDATA(index);

    wire [14:0] thalf_x0;
    wire [24:0] half_x03;
    assign thalf_x0 = tdata[39:25];
    assign half_x03 = tdata[24:0];

    wire [7:0] ey;
    assign ey = (ex == 0) ? 0: (8'd63 + {1'b0,ex[7:1]} + odd_flag - (x[23:3] == {1'b1,20'b0} & x[2:0] < 3'd6));

    // stage2
    wire [48:0] half_ax03;
    assign half_ax03 = {1'b1,mx_reg1} * half_x03_reg;

    // stage3
    wire [24:0] mra;
    assign mra = {thalf_x0_reg2,10'b0} - {1'b0,half_ax03_reg};

    wire [22:0] mr;
    assign mr = mra[22:0];

    // stage4
    wire [47:0] mya;
    assign mya = {1'b1,mr_reg} * {1'b1,mx_reg3};

    wire [22:0] my;
    assign my = (mya[47:47]) ? mya[46:24]: mya[45:23];

    always @(posedge clk) begin
        // stage1
        ey_reg1 <= ey;
        mx_reg1 <= mx;
        thalf_x0_reg1 <= thalf_x0;
        half_x03_reg <= half_x03;
        // stage2
        ey_reg2 <= ey_reg1;
        mx_reg2 <= mx_reg1;
        half_ax03_reg <= half_ax03[48:25];
        thalf_x0_reg2 <= thalf_x0_reg1;
        // stage3
        ey_reg3 <= ey_reg2;
        mx_reg3 <= mx_reg2;
        mr_reg <= mr;
        // stage4
        y <= {1'b0,ey_reg3,my};
    end

endmodule
