module finv(
    input wire [31:0] x,
    output wire [31:0] y
);

    function [36:0] TDATA (
	input [9:0] ML
    );
    begin
        casex(ML)
        10'd0: TDATA = 37'b1111111111000000000011111111111110000;
        10'd1: TDATA = 37'b1111111101000000010011111111111010000;
        10'd2: TDATA = 37'b1111111011000000110011111111110110000;
        10'd3: TDATA = 37'b1111111001000001100011011111110010000;
        10'd4: TDATA = 37'b1111110111000010100011011111101110000;
        10'd5: TDATA = 37'b1111110101000011110010011111101010000;
        10'd6: TDATA = 37'b1111110011000101010001111111100110001;
        10'd7: TDATA = 37'b1111110001000111000000011111100010001;
        10'd8: TDATA = 37'b1111101111001000111110111111011110100;
        10'd9: TDATA = 37'b1111101101001011001101011111011010100;
        10'd10: TDATA = 37'b1111101011001101101010111111010110100;
        10'd11: TDATA = 37'b1111101001010000011000011111010010111;
        10'd12: TDATA = 37'b1111100111010011010100111111001110111;
        10'd13: TDATA = 37'b1111100101010110100000111111001011000;
        10'd14: TDATA = 37'b1111100011011001111100011111000111001;
        10'd15: TDATA = 37'b1111100001011101100111011111000011011;
        10'd16: TDATA = 37'b1111011111100001100001011110111111100;
        10'd17: TDATA = 37'b1111011101100101101010111110111011101;
        10'd18: TDATA = 37'b1111011011101010000011011110111000000;
        10'd19: TDATA = 37'b1111011001101110101010111110110100000;
        10'd20: TDATA = 37'b1111010111110011100001111110110000011;
        10'd21: TDATA = 37'b1111010101111000100111111110101100100;
        10'd22: TDATA = 37'b1111010011111101111100111110101000111;
        10'd23: TDATA = 37'b1111010010000011100000111110100101000;
        10'd24: TDATA = 37'b1111010000001001010011111110100001011;
        10'd25: TDATA = 37'b1111001110001111010101011110011101100;
        10'd26: TDATA = 37'b1111001100010101100110011110011010000;
        10'd27: TDATA = 37'b1111001010011100000101111110010110011;
        10'd28: TDATA = 37'b1111001000100010110011111110010010100;
        10'd29: TDATA = 37'b1111000110101001110000111110001110111;
        10'd30: TDATA = 37'b1111000100110000111100111110001011001;
        10'd31: TDATA = 37'b1111000010111000010110111110000111100;
        10'd32: TDATA = 37'b1111000000111111111111111110000011111;
        10'd33: TDATA = 37'b1110111111000111110111011110000000001;
        10'd34: TDATA = 37'b1110111101001111111101011101111100100;
        10'd35: TDATA = 37'b1110111011011000010001111101111001000;
        10'd36: TDATA = 37'b1110111001100000110100111101110101100;
        10'd37: TDATA = 37'b1110110111101001100110011101110001111;
        10'd38: TDATA = 37'b1110110101110010100110011101101110001;
        10'd39: TDATA = 37'b1110110011111011110100011101101010100;
        10'd40: TDATA = 37'b1110110010000101010000111101100111000;
        10'd41: TDATA = 37'b1110110000001110111011011101100011100;
        10'd42: TDATA = 37'b1110101110011000110011111101100000000;
        10'd43: TDATA = 37'b1110101100100010111010111101011100100;
        10'd44: TDATA = 37'b1110101010101101001111111101011001000;
        10'd45: TDATA = 37'b1110101000110111110011011101010101011;
        10'd46: TDATA = 37'b1110100111000010100100011101010001111;
        10'd47: TDATA = 37'b1110100101001101100011111101001110100;
        10'd48: TDATA = 37'b1110100011011000110000111101001011000;
        10'd49: TDATA = 37'b1110100001100100001011111101000111100;
        10'd50: TDATA = 37'b1110011111101111110100111101000100000;
        10'd51: TDATA = 37'b1110011101111011101011111101000000100;
        10'd52: TDATA = 37'b1110011100000111110000011100111101000;
        10'd53: TDATA = 37'b1110011010010100000010111100111001101;
        10'd54: TDATA = 37'b1110011000100000100010111100110110001;
        10'd55: TDATA = 37'b1110010110101101010000111100110010111;
        10'd56: TDATA = 37'b1110010100111010001100011100101111011;
        10'd57: TDATA = 37'b1110010011000111010101011100101100000;
        10'd58: TDATA = 37'b1110010001010100101100011100101000100;
        10'd59: TDATA = 37'b1110001111100010010000011100100101001;
        10'd60: TDATA = 37'b1110001101110000000010011100100001111;
        10'd61: TDATA = 37'b1110001011111110000001011100011110100;
        10'd62: TDATA = 37'b1110001010001100001110011100011011001;
        10'd63: TDATA = 37'b1110001000011010101000011100010111101;
        10'd64: TDATA = 37'b1110000110101001001111111100010100100;
        10'd65: TDATA = 37'b1110000100111000000100011100010001001;
        10'd66: TDATA = 37'b1110000011000111000110011100001101101;
        10'd67: TDATA = 37'b1110000001010110010101111100001010100;
        10'd68: TDATA = 37'b1101111111100101110010011100000111001;
        10'd69: TDATA = 37'b1101111101110101011011111100000100000;
        10'd70: TDATA = 37'b1101111100000101010010111100000000100;
        10'd71: TDATA = 37'b1101111010010101010110011011111101011;
        10'd72: TDATA = 37'b1101111000100101100111011011111010000;
        10'd73: TDATA = 37'b1101110110110110000101011011110110111;
        10'd74: TDATA = 37'b1101110101000110110000011011110011100;
        10'd75: TDATA = 37'b1101110011010111101000011011110000011;
        10'd76: TDATA = 37'b1101110001101000101101011011101101001;
        10'd77: TDATA = 37'b1101101111111001111111011011101010000;
        10'd78: TDATA = 37'b1101101110001011011101111011100110101;
        10'd79: TDATA = 37'b1101101100011101001001011011100011100;
        10'd80: TDATA = 37'b1101101010101111000001011011100000011;
        10'd81: TDATA = 37'b1101101001000001000110011011011101001;
        10'd82: TDATA = 37'b1101100111010011010111111011011010000;
        10'd83: TDATA = 37'b1101100101100101110110011011010110111;
        10'd84: TDATA = 37'b1101100011111000100001011011010011101;
        10'd85: TDATA = 37'b1101100010001011011001011011010000100;
        10'd86: TDATA = 37'b1101100000011110011101011011001101011;
        10'd87: TDATA = 37'b1101011110110001101110011011001010001;
        10'd88: TDATA = 37'b1101011101000101001011011011000111000;
        10'd89: TDATA = 37'b1101011011011000110101011011000100000;
        10'd90: TDATA = 37'b1101011001101100101011011011000001000;
        10'd91: TDATA = 37'b1101011000000000101101111010111101111;
        10'd92: TDATA = 37'b1101010110010100111100111010111010101;
        10'd93: TDATA = 37'b1101010100101001011000011010110111100;
        10'd94: TDATA = 37'b1101010010111101111111111010110100100;
        10'd95: TDATA = 37'b1101010001010010110011111010110001100;
        10'd96: TDATA = 37'b1101001111100111110011111010101110011;
        10'd97: TDATA = 37'b1101001101111101000000011010101011011;
        10'd98: TDATA = 37'b1101001100010010011000111010101000011;
        10'd99: TDATA = 37'b1101001010100111111101011010100101001;
        10'd100: TDATA = 37'b1101001000111101101110011010100010001;
        10'd101: TDATA = 37'b1101000111010011101011011010011111001;
        10'd102: TDATA = 37'b1101000101101001110100011010011100001;
        10'd103: TDATA = 37'b1101000100000000001001011010011001011;
        10'd104: TDATA = 37'b1101000010010110101001111010010110001;
        10'd105: TDATA = 37'b1101000000101101010110111010010011001;
        10'd106: TDATA = 37'b1100111111000100001111111010010000011;
        10'd107: TDATA = 37'b1100111101011011010100011010001101001;
        10'd108: TDATA = 37'b1100111011110010100100111010001010011;
        10'd109: TDATA = 37'b1100111010001010000001011010000111011;
        10'd110: TDATA = 37'b1100111000100001101001111010000100100;
        10'd111: TDATA = 37'b1100110110111001011101111010000001100;
        10'd112: TDATA = 37'b1100110101010001011101011001111110100;
        10'd113: TDATA = 37'b1100110011101001101000111001111011101;
        10'd114: TDATA = 37'b1100110010000001111111111001111000101;
        10'd115: TDATA = 37'b1100110000011010100010011001110101111;
        10'd116: TDATA = 37'b1100101110110011010000111001110011000;
        10'd117: TDATA = 37'b1100101101001100001010111001110000000;
        10'd118: TDATA = 37'b1100101011100101010000011001101101001;
        10'd119: TDATA = 37'b1100101001111110100001011001101010001;
        10'd120: TDATA = 37'b1100101000010111111101111001100111011;
        10'd121: TDATA = 37'b1100100110110001100101011001100100100;
        10'd122: TDATA = 37'b1100100101001011011000111001100001101;
        10'd123: TDATA = 37'b1100100011100101010111111001011110111;
        10'd124: TDATA = 37'b1100100001111111100001111001011100000;
        10'd125: TDATA = 37'b1100100000011001110111011001011001001;
        10'd126: TDATA = 37'b1100011110110100010111111001010110100;
        10'd127: TDATA = 37'b1100011101001111000011111001010011100;
        10'd128: TDATA = 37'b1100011011101001111011011001010000101;
        10'd129: TDATA = 37'b1100011010000100111101111001001110000;
        10'd130: TDATA = 37'b1100011000100000001011111001001011001;
        10'd131: TDATA = 37'b1100010110111011100100011001001000011;
        10'd132: TDATA = 37'b1100010101010111001000011001000101100;
        10'd133: TDATA = 37'b1100010011110010110111111001000010111;
        10'd134: TDATA = 37'b1100010010001110110001111001000000000;
        10'd135: TDATA = 37'b1100010000101010110111011000111101001;
        10'd136: TDATA = 37'b1100001111000111000111011000111010100;
        10'd137: TDATA = 37'b1100001101100011100010111000110111101;
        10'd138: TDATA = 37'b1100001100000000001000111000110101000;
        10'd139: TDATA = 37'b1100001010011100111001111000110010011;
        10'd140: TDATA = 37'b1100001000111001110110011000101111100;
        10'd141: TDATA = 37'b1100000111010110111101011000101100111;
        10'd142: TDATA = 37'b1100000101110100001110111000101010001;
        10'd143: TDATA = 37'b1100000100010001101011011000100111100;
        10'd144: TDATA = 37'b1100000010101111010010111000100100101;
        10'd145: TDATA = 37'b1100000001001101000101011000100010000;
        10'd146: TDATA = 37'b1011111111101011000001111000011111011;
        10'd147: TDATA = 37'b1011111110001001001001111000011100101;
        10'd148: TDATA = 37'b1011111100100111011011111000011010000;
        10'd149: TDATA = 37'b1011111011000101111000111000010111011;
        10'd150: TDATA = 37'b1011111001100100100000111000010100111;
        10'd151: TDATA = 37'b1011111000000011010010111000010010000;
        10'd152: TDATA = 37'b1011110110100010001111111000001111100;
        10'd153: TDATA = 37'b1011110101000001010110111000001100111;
        10'd154: TDATA = 37'b1011110011100000101000111000001010001;
        10'd155: TDATA = 37'b1011110010000000000101011000000111100;
        10'd156: TDATA = 37'b1011110000011111101100011000000101000;
        10'd157: TDATA = 37'b1011101110111111011101011000000010011;
        10'd158: TDATA = 37'b1011101101011111011001010111111111101;
        10'd159: TDATA = 37'b1011101011111111011111010111111101000;
        10'd160: TDATA = 37'b1011101010011111101111110111111010100;
        10'd161: TDATA = 37'b1011101001000000001010010111111000000;
        10'd162: TDATA = 37'b1011100111100000101111010111110101100;
        10'd163: TDATA = 37'b1011100110000001011110110111110010111;
        10'd164: TDATA = 37'b1011100100100010011000110111110000001;
        10'd165: TDATA = 37'b1011100011000011011100010111101101101;
        10'd166: TDATA = 37'b1011100001100100101010010111101011001;
        10'd167: TDATA = 37'b1011100000000110000010110111101000100;
        10'd168: TDATA = 37'b1011011110100111100101010111100110000;
        10'd169: TDATA = 37'b1011011101001001010001110111100011100;
        10'd170: TDATA = 37'b1011011011101011001000010111100001000;
        10'd171: TDATA = 37'b1011011010001101001001010111011110100;
        10'd172: TDATA = 37'b1011011000101111010011110111011100000;
        10'd173: TDATA = 37'b1011010111010001101000110111011001100;
        10'd174: TDATA = 37'b1011010101110100000111110111010111000;
        10'd175: TDATA = 37'b1011010100010110110000010111010100100;
        10'd176: TDATA = 37'b1011010010111001100011010111010010000;
        10'd177: TDATA = 37'b1011010001011100011111110111001111100;
        10'd178: TDATA = 37'b1011001111111111100110110111001101000;
        10'd179: TDATA = 37'b1011001110100010110110110111001010100;
        10'd180: TDATA = 37'b1011001101000110010001010111001000001;
        10'd181: TDATA = 37'b1011001011101001110101010111000101101;
        10'd182: TDATA = 37'b1011001010001101100011010111000011001;
        10'd183: TDATA = 37'b1011001000110001011011010111000000111;
        10'd184: TDATA = 37'b1011000111010101011100110110111110011;
        10'd185: TDATA = 37'b1011000101111001100111110110111100000;
        10'd186: TDATA = 37'b1011000100011101111100110110111001100;
        10'd187: TDATA = 37'b1011000011000010011011110110110111000;
        10'd188: TDATA = 37'b1011000001100111000011110110110100101;
        10'd189: TDATA = 37'b1011000000001011110101110110110010001;
        10'd190: TDATA = 37'b1010111110110000110001010110110000000;
        10'd191: TDATA = 37'b1010111101010101110110110110101101100;
        10'd192: TDATA = 37'b1010111011111011000101010110101011000;
        10'd193: TDATA = 37'b1010111010100000011101110110101000101;
        10'd194: TDATA = 37'b1010111001000101111111010110100110011;
        10'd195: TDATA = 37'b1010110111101011101010110110100100000;
        10'd196: TDATA = 37'b1010110110010001011111010110100001100;
        10'd197: TDATA = 37'b1010110100110111011101010110011111001;
        10'd198: TDATA = 37'b1010110011011101100101010110011101000;
        10'd199: TDATA = 37'b1010110010000011110110010110011010100;
        10'd200: TDATA = 37'b1010110000101010010000110110011000001;
        10'd201: TDATA = 37'b1010101111010000110100010110010101111;
        10'd202: TDATA = 37'b1010101101110111100001010110010011100;
        10'd203: TDATA = 37'b1010101100011110010111110110010001001;
        10'd204: TDATA = 37'b1010101011000101010111110110001111000;
        10'd205: TDATA = 37'b1010101001101100100000010110001100100;
        10'd206: TDATA = 37'b1010101000010011110010110110001010001;
        10'd207: TDATA = 37'b1010100110111011001110010110001000000;
        10'd208: TDATA = 37'b1010100101100010110010110110000101100;
        10'd209: TDATA = 37'b1010100100001010100000110110000011011;
        10'd210: TDATA = 37'b1010100010110010010111010110000001000;
        10'd211: TDATA = 37'b1010100001011010010111110101111110111;
        10'd212: TDATA = 37'b1010100000000010100000110101111100100;
        10'd213: TDATA = 37'b1010011110101010110011010101111010001;
        10'd214: TDATA = 37'b1010011101010011001110010101111000000;
        10'd215: TDATA = 37'b1010011011111011110010110101110101101;
        10'd216: TDATA = 37'b1010011010100100100000010101110011100;
        10'd217: TDATA = 37'b1010011001001101010110110101110001001;
        10'd218: TDATA = 37'b1010010111110110010101110101101111000;
        10'd219: TDATA = 37'b1010010110011111011110010101101100101;
        10'd220: TDATA = 37'b1010010101001000101111110101101010100;
        10'd221: TDATA = 37'b1010010011110010001001110101101000011;
        10'd222: TDATA = 37'b1010010010011011101100110101100110000;
        10'd223: TDATA = 37'b1010010001000101011000110101100011111;
        10'd224: TDATA = 37'b1010001111101111001101110101100001100;
        10'd225: TDATA = 37'b1010001110011001001011010101011111100;
        10'd226: TDATA = 37'b1010001101000011010001110101011101001;
        10'd227: TDATA = 37'b1010001011101101100000110101011011000;
        10'd228: TDATA = 37'b1010001010010111111000110101011000111;
        10'd229: TDATA = 37'b1010001001000010011001110101010110101;
        10'd230: TDATA = 37'b1010000111101101000011010101010100100;
        10'd231: TDATA = 37'b1010000110010111110101010101010010011;
        10'd232: TDATA = 37'b1010000101000010110000010101010000001;
        10'd233: TDATA = 37'b1010000011101101110011110101001110000;
        10'd234: TDATA = 37'b1010000010011000111111110101001011111;
        10'd235: TDATA = 37'b1010000001000100010100110101001001101;
        10'd236: TDATA = 37'b1001111111101111110001110101000111100;
        10'd237: TDATA = 37'b1001111110011011010111110101000101011;
        10'd238: TDATA = 37'b1001111101000111000110010101000011001;
        10'd239: TDATA = 37'b1001111011110010111101010101000001000;
        10'd240: TDATA = 37'b1001111010011110111100110100111111000;
        10'd241: TDATA = 37'b1001111001001011000100110100111100111;
        10'd242: TDATA = 37'b1001110111110111010101010100111010101;
        10'd243: TDATA = 37'b1001110110100011101110010100111000100;
        10'd244: TDATA = 37'b1001110101010000001111110100110110100;
        10'd245: TDATA = 37'b1001110011111100111001110100110100100;
        10'd246: TDATA = 37'b1001110010101001101011110100110010011;
        10'd247: TDATA = 37'b1001110001010110100110110100110000001;
        10'd248: TDATA = 37'b1001110000000011101001110100101110001;
        10'd249: TDATA = 37'b1001101110110000110100110100101100000;
        10'd250: TDATA = 37'b1001101101011110001000010100101010000;
        10'd251: TDATA = 37'b1001101100001011100100010100101000000;
        10'd252: TDATA = 37'b1001101010111001001000110100100110000;
        10'd253: TDATA = 37'b1001101001100110110101010100100011111;
        10'd254: TDATA = 37'b1001101000010100101001110100100001111;
        10'd255: TDATA = 37'b1001100111000010100110110100011111101;
        10'd256: TDATA = 37'b1001100101110000101011110100011101101;
        10'd257: TDATA = 37'b1001100100011110111001010100011011100;
        10'd258: TDATA = 37'b1001100011001101001110110100011001100;
        10'd259: TDATA = 37'b1001100001111011101100010100010111100;
        10'd260: TDATA = 37'b1001100000101010010001110100010101100;
        10'd261: TDATA = 37'b1001011111011000111111110100010011100;
        10'd262: TDATA = 37'b1001011110000111110101110100010001100;
        10'd263: TDATA = 37'b1001011100110110110011110100001111100;
        10'd264: TDATA = 37'b1001011011100101111001110100001101100;
        10'd265: TDATA = 37'b1001011010010101000111110100001011100;
        10'd266: TDATA = 37'b1001011001000100011101110100001001100;
        10'd267: TDATA = 37'b1001010111110011111011110100000111100;
        10'd268: TDATA = 37'b1001010110100011100001110100000101100;
        10'd269: TDATA = 37'b1001010101010011001111110100000011100;
        10'd270: TDATA = 37'b1001010100000011000101110100000001100;
        10'd271: TDATA = 37'b1001010010110011000011110011111111100;
        10'd272: TDATA = 37'b1001010001100011001001110011111101100;
        10'd273: TDATA = 37'b1001010000010011010111010011111011100;
        10'd274: TDATA = 37'b1001001111000011101100110011111001100;
        10'd275: TDATA = 37'b1001001101110100001010010011110111101;
        10'd276: TDATA = 37'b1001001100100100101111010011110101101;
        10'd277: TDATA = 37'b1001001011010101011100010011110011101;
        10'd278: TDATA = 37'b1001001010000110010001010011110001111;
        10'd279: TDATA = 37'b1001001000110111001101110011101111111;
        10'd280: TDATA = 37'b1001000111101000010010010011101110000;
        10'd281: TDATA = 37'b1001000110011001011110010011101100000;
        10'd282: TDATA = 37'b1001000101001010110001110011101010000;
        10'd283: TDATA = 37'b1001000011111100001101010011101000001;
        10'd284: TDATA = 37'b1001000010101101110000110011100110001;
        10'd285: TDATA = 37'b1001000001011111011011010011100100001;
        10'd286: TDATA = 37'b1001000000010001001101110011100010100;
        10'd287: TDATA = 37'b1000111111000011001000010011100000100;
        10'd288: TDATA = 37'b1000111101110101001001110011011110100;
        10'd289: TDATA = 37'b1000111100100111010011010011011100101;
        10'd290: TDATA = 37'b1000111011011001100100010011011010111;
        10'd291: TDATA = 37'b1000111010001011111100110011011000111;
        10'd292: TDATA = 37'b1000111000111110011100110011010111000;
        10'd293: TDATA = 37'b1000110111110001000100010011010101001;
        10'd294: TDATA = 37'b1000110110100011110011010011010011001;
        10'd295: TDATA = 37'b1000110101010110101001110011010001011;
        10'd296: TDATA = 37'b1000110100001001100111110011001111100;
        10'd297: TDATA = 37'b1000110010111100101101010011001101101;
        10'd298: TDATA = 37'b1000110001101111111010010011001011101;
        10'd299: TDATA = 37'b1000110000100011001110110011001010000;
        10'd300: TDATA = 37'b1000101111010110101010110011001000000;
        10'd301: TDATA = 37'b1000101110001010001101110011000110001;
        10'd302: TDATA = 37'b1000101100111101111000010011000100100;
        10'd303: TDATA = 37'b1000101011110001101010010011000010100;
        10'd304: TDATA = 37'b1000101010100101100011110011000000101;
        10'd305: TDATA = 37'b1000101001011001100100010010111111000;
        10'd306: TDATA = 37'b1000101000001101101100010010111101000;
        10'd307: TDATA = 37'b1000100111000001111011010010111011001;
        10'd308: TDATA = 37'b1000100101110110010001110010111001100;
        10'd309: TDATA = 37'b1000100100101010101111010010110111100;
        10'd310: TDATA = 37'b1000100011011111010100010010110101111;
        10'd311: TDATA = 37'b1000100010010100000000110010110100000;
        10'd312: TDATA = 37'b1000100001001000110100010010110010001;
        10'd313: TDATA = 37'b1000011111111101101110110010110000100;
        10'd314: TDATA = 37'b1000011110110010110000110010101110100;
        10'd315: TDATA = 37'b1000011101100111111001110010101100111;
        10'd316: TDATA = 37'b1000011100011101001001110010101011000;
        10'd317: TDATA = 37'b1000011011010010100000110010101001001;
        10'd318: TDATA = 37'b1000011010000111111111010010100111100;
        10'd319: TDATA = 37'b1000011000111101100100110010100101101;
        10'd320: TDATA = 37'b1000010111110011010001010010100100000;
        10'd321: TDATA = 37'b1000010110101001000100110010100010001;
        10'd322: TDATA = 37'b1000010101011110111111110010100000100;
        10'd323: TDATA = 37'b1000010100010101000001010010011110101;
        10'd324: TDATA = 37'b1000010011001011001010010010011100111;
        10'd325: TDATA = 37'b1000010010000001011001110010011011001;
        10'd326: TDATA = 37'b1000010000110111110000110010011001011;
        10'd327: TDATA = 37'b1000001111101110001110010010010111101;
        10'd328: TDATA = 37'b1000001110100100110010110010010110000;
        10'd329: TDATA = 37'b1000001101011011011110010010010100001;
        10'd330: TDATA = 37'b1000001100010010010001010010010010100;
        10'd331: TDATA = 37'b1000001011001001001010010010010000101;
        10'd332: TDATA = 37'b1000001010000000001010110010001111000;
        10'd333: TDATA = 37'b1000001000110111010010010010001101011;
        10'd334: TDATA = 37'b1000000111101110100000010010001011100;
        10'd335: TDATA = 37'b1000000110100101110101010010001001111;
        10'd336: TDATA = 37'b1000000101011101010000110010001000001;
        10'd337: TDATA = 37'b1000000100010100110011010010000110100;
        10'd338: TDATA = 37'b1000000011001100011100110010000100111;
        10'd339: TDATA = 37'b1000000010000100001101010010000011000;
        10'd340: TDATA = 37'b1000000000111100000100010010000001100;
        10'd341: TDATA = 37'b0111111111110100000001110001111111101;
        10'd342: TDATA = 37'b0111111110101100000110010001111110000;
        10'd343: TDATA = 37'b0111111101100100010001110001111100011;
        10'd344: TDATA = 37'b0111111100011100100011110001111010101;
        10'd345: TDATA = 37'b0111111011010100111100010001111001000;
        10'd346: TDATA = 37'b0111111010001101011011110001110111011;
        10'd347: TDATA = 37'b0111111001000110000001110001110101100;
        10'd348: TDATA = 37'b0111110111111110101110010001110100000;
        10'd349: TDATA = 37'b0111110110110111100001110001110010011;
        10'd350: TDATA = 37'b0111110101110000011011010001110000101;
        10'd351: TDATA = 37'b0111110100101001011100010001101111000;
        10'd352: TDATA = 37'b0111110011100010100011010001101101011;
        10'd353: TDATA = 37'b0111110010011011110000110001101011101;
        10'd354: TDATA = 37'b0111110001010101000101010001101010000;
        10'd355: TDATA = 37'b0111110000001110100000010001101000100;
        10'd356: TDATA = 37'b0111101111001000000001110001100110111;
        10'd357: TDATA = 37'b0111101110000001101001110001100101001;
        10'd358: TDATA = 37'b0111101100111011010111110001100011100;
        10'd359: TDATA = 37'b0111101011110101001100110001100010000;
        10'd360: TDATA = 37'b0111101010101111001000010001100000011;
        10'd361: TDATA = 37'b0111101001101001001010010001011110101;
        10'd362: TDATA = 37'b0111101000100011010010110001011101000;
        10'd363: TDATA = 37'b0111100111011101100001110001011011100;
        10'd364: TDATA = 37'b0111100110010111110110110001011001111;
        10'd365: TDATA = 37'b0111100101010010010010110001011000001;
        10'd366: TDATA = 37'b0111100100001100110100110001010110101;
        10'd367: TDATA = 37'b0111100011000111011101010001010101000;
        10'd368: TDATA = 37'b0111100010000010001011110001010011100;
        10'd369: TDATA = 37'b0111100000111101000001010001010010000;
        10'd370: TDATA = 37'b0111011111110111111100110001010000001;
        10'd371: TDATA = 37'b0111011110110010111110110001001110101;
        10'd372: TDATA = 37'b0111011101101110000110110001001101000;
        10'd373: TDATA = 37'b0111011100101001010101010001001011100;
        10'd374: TDATA = 37'b0111011011100100101010010001001010000;
        10'd375: TDATA = 37'b0111011010100000000101010001001000100;
        10'd376: TDATA = 37'b0111011001011011100110110001000110111;
        10'd377: TDATA = 37'b0111011000010111001110010001000101001;
        10'd378: TDATA = 37'b0111010111010010111100010001000011101;
        10'd379: TDATA = 37'b0111010110001110110000010001000010001;
        10'd380: TDATA = 37'b0111010101001010101010110001000000100;
        10'd381: TDATA = 37'b0111010100000110101011010000111111000;
        10'd382: TDATA = 37'b0111010011000010110001110000111101100;
        10'd383: TDATA = 37'b0111010001111110111110110000111100000;
        10'd384: TDATA = 37'b0111010000111011010001110000111010100;
        10'd385: TDATA = 37'b0111001111110111101011010000111000111;
        10'd386: TDATA = 37'b0111001110110100001010010000110111100;
        10'd387: TDATA = 37'b0111001101110000101111110000110101111;
        10'd388: TDATA = 37'b0111001100101101011011010000110100011;
        10'd389: TDATA = 37'b0111001011101010001101010000110010111;
        10'd390: TDATA = 37'b0111001010100111000100110000110001001;
        10'd391: TDATA = 37'b0111001001100100000010110000101111111;
        10'd392: TDATA = 37'b0111001000100001000110010000101110011;
        10'd393: TDATA = 37'b0111000111011110010000010000101100101;
        10'd394: TDATA = 37'b0111000110011011100000010000101011001;
        10'd395: TDATA = 37'b0111000101011000110110010000101001101;
        10'd396: TDATA = 37'b0111000100010110010010010000101000001;
        10'd397: TDATA = 37'b0111000011010011110100010000100110101;
        10'd398: TDATA = 37'b0111000010010001011100010000100101001;
        10'd399: TDATA = 37'b0111000001001111001010010000100011101;
        10'd400: TDATA = 37'b0111000000001100111101110000100010011;
        10'd401: TDATA = 37'b0110111111001010110111110000100000101;
        10'd402: TDATA = 37'b0110111110001000110111010000011111011;
        10'd403: TDATA = 37'b0110111101000110111101010000011101111;
        10'd404: TDATA = 37'b0110111100000101001000110000011100011;
        10'd405: TDATA = 37'b0110111011000011011010010000011010111;
        10'd406: TDATA = 37'b0110111010000001110001010000011001100;
        10'd407: TDATA = 37'b0110111001000000001110110000011000000;
        10'd408: TDATA = 37'b0110110111111110110001110000010110100;
        10'd409: TDATA = 37'b0110110110111101011010110000010101000;
        10'd410: TDATA = 37'b0110110101111100001001010000010011100;
        10'd411: TDATA = 37'b0110110100111010111101110000010010000;
        10'd412: TDATA = 37'b0110110011111001111000010000010000101;
        10'd413: TDATA = 37'b0110110010111000111000010000001111001;
        10'd414: TDATA = 37'b0110110001110111111110010000001101101;
        10'd415: TDATA = 37'b0110110000110111001010010000001100011;
        10'd416: TDATA = 37'b0110101111110110011011110000001010111;
        10'd417: TDATA = 37'b0110101110110101110010110000001001100;
        10'd418: TDATA = 37'b0110101101110101001111110000001000000;
        10'd419: TDATA = 37'b0110101100110100110010010000000110100;
        10'd420: TDATA = 37'b0110101011110100011010110000000101001;
        10'd421: TDATA = 37'b0110101010110100001000110000000011111;
        10'd422: TDATA = 37'b0110101001110011111100110000000010011;
        10'd423: TDATA = 37'b0110101000110011110110010000000000111;
        10'd424: TDATA = 37'b0110100111110011110101001111111111100;
        10'd425: TDATA = 37'b0110100110110011111010001111111110000;
        10'd426: TDATA = 37'b0110100101110100000100001111111100101;
        10'd427: TDATA = 37'b0110100100110100010100101111111011011;
        10'd428: TDATA = 37'b0110100011110100101010001111111001111;
        10'd429: TDATA = 37'b0110100010110101000101001111111000100;
        10'd430: TDATA = 37'b0110100001110101100110001111110111000;
        10'd431: TDATA = 37'b0110100000110110001100101111110101101;
        10'd432: TDATA = 37'b0110011111110110111000101111110100001;
        10'd433: TDATA = 37'b0110011110110111101010001111110010111;
        10'd434: TDATA = 37'b0110011101111000100001101111110001100;
        10'd435: TDATA = 37'b0110011100111001011110001111110000000;
        10'd436: TDATA = 37'b0110011011111010100000001111101110101;
        10'd437: TDATA = 37'b0110011010111011101000001111101101011;
        10'd438: TDATA = 37'b0110011001111100110101001111101100000;
        10'd439: TDATA = 37'b0110011000111110001000001111101010100;
        10'd440: TDATA = 37'b0110010111111111100000001111101001001;
        10'd441: TDATA = 37'b0110010111000000111101101111101000000;
        10'd442: TDATA = 37'b0110010110000010100000101111100110100;
        10'd443: TDATA = 37'b0110010101000100001001101111100101001;
        10'd444: TDATA = 37'b0110010100000101110111101111100011111;
        10'd445: TDATA = 37'b0110010011000111101010101111100010100;
        10'd446: TDATA = 37'b0110010010001001100011101111100001000;
        10'd447: TDATA = 37'b0110010001001011100010001111011111101;
        10'd448: TDATA = 37'b0110010000001101100101101111011110100;
        10'd449: TDATA = 37'b0110001111001111101110101111011101000;
        10'd450: TDATA = 37'b0110001110010001111101001111011011101;
        10'd451: TDATA = 37'b0110001101010100010000101111011010100;
        10'd452: TDATA = 37'b0110001100010110101001101111011001000;
        10'd453: TDATA = 37'b0110001011011001001000001111010111101;
        10'd454: TDATA = 37'b0110001010011011101100001111010110011;
        10'd455: TDATA = 37'b0110001001011110010101001111010101000;
        10'd456: TDATA = 37'b0110001000100001000011001111010011101;
        10'd457: TDATA = 37'b0110000111100011110111001111010010011;
        10'd458: TDATA = 37'b0110000110100110110000001111010001000;
        10'd459: TDATA = 37'b0110000101101001101110001111001111101;
        10'd460: TDATA = 37'b0110000100101100110001101111001110100;
        10'd461: TDATA = 37'b0110000011101111111010101111001101000;
        10'd462: TDATA = 37'b0110000010110011001000001111001011111;
        10'd463: TDATA = 37'b0110000001110110011011101111001010100;
        10'd464: TDATA = 37'b0110000000111001110100001111001001001;
        10'd465: TDATA = 37'b0101111111111101010001101111001000000;
        10'd466: TDATA = 37'b0101111111000000110100101111000110101;
        10'd467: TDATA = 37'b0101111110000100011100101111000101011;
        10'd468: TDATA = 37'b0101111101001000001001101111000100000;
        10'd469: TDATA = 37'b0101111100001011111100001111000010101;
        10'd470: TDATA = 37'b0101111011001111110011101111000001100;
        10'd471: TDATA = 37'b0101111010010011110000001111000000000;
        10'd472: TDATA = 37'b0101111001010111110010001110111110111;
        10'd473: TDATA = 37'b0101111000011011111001001110111101100;
        10'd474: TDATA = 37'b0101110111100000000101001110111100011;
        10'd475: TDATA = 37'b0101110110100100010110001110111011000;
        10'd476: TDATA = 37'b0101110101101000101100101110111001111;
        10'd477: TDATA = 37'b0101110100101101000111101110111000100;
        10'd478: TDATA = 37'b0101110011110001101000001110110111001;
        10'd479: TDATA = 37'b0101110010110110001101101110110110000;
        10'd480: TDATA = 37'b0101110001111010111000001110110100101;
        10'd481: TDATA = 37'b0101110000111111100111101110110011100;
        10'd482: TDATA = 37'b0101110000000100011100101110110010001;
        10'd483: TDATA = 37'b0101101111001001010110001110110001000;
        10'd484: TDATA = 37'b0101101110001110010100101110101111101;
        10'd485: TDATA = 37'b0101101101010011011000001110101110100;
        10'd486: TDATA = 37'b0101101100011000100001001110101101001;
        10'd487: TDATA = 37'b0101101011011101101110101110101100000;
        10'd488: TDATA = 37'b0101101010100011000001001110101010101;
        10'd489: TDATA = 37'b0101101001101000011000101110101001100;
        10'd490: TDATA = 37'b0101101000101101110101001110101000001;
        10'd491: TDATA = 37'b0101100111110011010110101110100111000;
        10'd492: TDATA = 37'b0101100110111000111101001110100101111;
        10'd493: TDATA = 37'b0101100101111110101000101110100100100;
        10'd494: TDATA = 37'b0101100101000100011000101110100011011;
        10'd495: TDATA = 37'b0101100100001010001110001110100010000;
        10'd496: TDATA = 37'b0101100011010000001000001110100000111;
        10'd497: TDATA = 37'b0101100010010110000111001110011111100;
        10'd498: TDATA = 37'b0101100001011100001010101110011110100;
        10'd499: TDATA = 37'b0101100000100010010011101110011101001;
        10'd500: TDATA = 37'b0101011111101000100001001110011100000;
        10'd501: TDATA = 37'b0101011110101110110011101110011010101;
        10'd502: TDATA = 37'b0101011101110101001010101110011001100;
        10'd503: TDATA = 37'b0101011100111011100110101110011000011;
        10'd504: TDATA = 37'b0101011100000010000111101110010111001;
        10'd505: TDATA = 37'b0101011011001000101101001110010110000;
        10'd506: TDATA = 37'b0101011010001111010111101110010100101;
        10'd507: TDATA = 37'b0101011001010110000111001110010011100;
        10'd508: TDATA = 37'b0101011000011100111011001110010010011;
        10'd509: TDATA = 37'b0101010111100011110100001110010001000;
        10'd510: TDATA = 37'b0101010110101010110001101110010000000;
        10'd511: TDATA = 37'b0101010101110001110100001110001110111;
        10'd512: TDATA = 37'b0101010100111000111011001110001101100;
        10'd513: TDATA = 37'b0101010100000000000111001110001100100;
        10'd514: TDATA = 37'b0101010011000111010111101110001011001;
        10'd515: TDATA = 37'b0101010010001110101100101110001010000;
        10'd516: TDATA = 37'b0101010001010110000110101110001000111;
        10'd517: TDATA = 37'b0101010000011101100101101110000111101;
        10'd518: TDATA = 37'b0101001111100101001001001110000110100;
        10'd519: TDATA = 37'b0101001110101100110001001110000101100;
        10'd520: TDATA = 37'b0101001101110100011101101110000100001;
        10'd521: TDATA = 37'b0101001100111100001111001110000011000;
        10'd522: TDATA = 37'b0101001100000100000101001110000010000;
        10'd523: TDATA = 37'b0101001011001100000000001110000000101;
        10'd524: TDATA = 37'b0101001010010011111111001101111111100;
        10'd525: TDATA = 37'b0101001001011100000011001101111110100;
        10'd526: TDATA = 37'b0101001000100100001011101101111101011;
        10'd527: TDATA = 37'b0101000111101100011001001101111100000;
        10'd528: TDATA = 37'b0101000110110100101010101101111011000;
        10'd529: TDATA = 37'b0101000101111101000001001101111001111;
        10'd530: TDATA = 37'b0101000101000101011100001101111000101;
        10'd531: TDATA = 37'b0101000100001101111011101101110111100;
        10'd532: TDATA = 37'b0101000011010110011111101101110110011;
        10'd533: TDATA = 37'b0101000010011111001000101101110101001;
        10'd534: TDATA = 37'b0101000001100111110101101101110100000;
        10'd535: TDATA = 37'b0101000000110000100111101101110011000;
        10'd536: TDATA = 37'b0100111111111001011101101101110001111;
        10'd537: TDATA = 37'b0100111111000010011000101101110000101;
        10'd538: TDATA = 37'b0100111110001011010111101101101111100;
        10'd539: TDATA = 37'b0100111101010100011011101101101110100;
        10'd540: TDATA = 37'b0100111100011101100100001101101101011;
        10'd541: TDATA = 37'b0100111011100110110000101101101100001;
        10'd542: TDATA = 37'b0100111010110000000010001101101011000;
        10'd543: TDATA = 37'b0100111001111001010111101101101010000;
        10'd544: TDATA = 37'b0100111001000010110010001101101000111;
        10'd545: TDATA = 37'b0100111000001100010000101101100111111;
        10'd546: TDATA = 37'b0100110111010101110011101101100110101;
        10'd547: TDATA = 37'b0100110110011111011011001101100101100;
        10'd548: TDATA = 37'b0100110101101001000111001101100100100;
        10'd549: TDATA = 37'b0100110100110010110111101101100011011;
        10'd550: TDATA = 37'b0100110011111100101100001101100010001;
        10'd551: TDATA = 37'b0100110011000110100101101101100001000;
        10'd552: TDATA = 37'b0100110010010000100011001101100000000;
        10'd553: TDATA = 37'b0100110001011010100101001101011111000;
        10'd554: TDATA = 37'b0100110000100100101011101101011101111;
        10'd555: TDATA = 37'b0100101111101110110110001101011100101;
        10'd556: TDATA = 37'b0100101110111001000101001101011011101;
        10'd557: TDATA = 37'b0100101110000011011000101101011010100;
        10'd558: TDATA = 37'b0100101101001101110000001101011001100;
        10'd559: TDATA = 37'b0100101100011000001100101101011000100;
        10'd560: TDATA = 37'b0100101011100010101101001101010111011;
        10'd561: TDATA = 37'b0100101010101101010001101101010110001;
        10'd562: TDATA = 37'b0100101001110111111010101101010101000;
        10'd563: TDATA = 37'b0100101001000010101000001101010100000;
        10'd564: TDATA = 37'b0100101000001101011001101101010011000;
        10'd565: TDATA = 37'b0100100111011000001111101101010010000;
        10'd566: TDATA = 37'b0100100110100011001001101101010000111;
        10'd567: TDATA = 37'b0100100101101110001000001101001111111;
        10'd568: TDATA = 37'b0100100100111001001011001101001110111;
        10'd569: TDATA = 37'b0100100100000100010010001101001101101;
        10'd570: TDATA = 37'b0100100011001111011101001101001100100;
        10'd571: TDATA = 37'b0100100010011010101100101101001011100;
        10'd572: TDATA = 37'b0100100001100110000000101101001010100;
        10'd573: TDATA = 37'b0100100000110001011000101101001001100;
        10'd574: TDATA = 37'b0100011111111100110100101101001000100;
        10'd575: TDATA = 37'b0100011111001000010101001101000111100;
        10'd576: TDATA = 37'b0100011110010011111001101101000110011;
        10'd577: TDATA = 37'b0100011101011111100010001101000101001;
        10'd578: TDATA = 37'b0100011100101011001111001101000100001;
        10'd579: TDATA = 37'b0100011011110111000000001101000011001;
        10'd580: TDATA = 37'b0100011011000010110101101101000010000;
        10'd581: TDATA = 37'b0100011010001110101111001101000001000;
        10'd582: TDATA = 37'b0100011001011010101100101101000000000;
        10'd583: TDATA = 37'b0100011000100110101110001100111111000;
        10'd584: TDATA = 37'b0100010111110010110100001100111110000;
        10'd585: TDATA = 37'b0100010110111110111110001100111101000;
        10'd586: TDATA = 37'b0100010110001011001100001100111100000;
        10'd587: TDATA = 37'b0100010101010111011110101100111010111;
        10'd588: TDATA = 37'b0100010100100011110100101100111001111;
        10'd589: TDATA = 37'b0100010011110000001111001100111001000;
        10'd590: TDATA = 37'b0100010010111100101101101100110111111;
        10'd591: TDATA = 37'b0100010010001001010000101100110110111;
        10'd592: TDATA = 37'b0100010001010101110111001100110101111;
        10'd593: TDATA = 37'b0100010000100010100001101100110100111;
        10'd594: TDATA = 37'b0100001111101111010000101100110011101;
        10'd595: TDATA = 37'b0100001110111100000011101100110010111;
        10'd596: TDATA = 37'b0100001110001000111010001100110001111;
        10'd597: TDATA = 37'b0100001101010101110101001100110000101;
        10'd598: TDATA = 37'b0100001100100010110100001100101111101;
        10'd599: TDATA = 37'b0100001011101111110111001100101110101;
        10'd600: TDATA = 37'b0100001010111100111110001100101101101;
        10'd601: TDATA = 37'b0100001010001010001001001100101100101;
        10'd602: TDATA = 37'b0100001001010111011000001100101011101;
        10'd603: TDATA = 37'b0100001000100100101011001100101010101;
        10'd604: TDATA = 37'b0100000111110010000010001100101001101;
        10'd605: TDATA = 37'b0100000110111111011101001100101000101;
        10'd606: TDATA = 37'b0100000110001100111100001100100111111;
        10'd607: TDATA = 37'b0100000101011010011111001100100110101;
        10'd608: TDATA = 37'b0100000100101000000101101100100101111;
        10'd609: TDATA = 37'b0100000011110101110000101100100100111;
        10'd610: TDATA = 37'b0100000011000011011111101100100011111;
        10'd611: TDATA = 37'b0100000010010001010010001100100010111;
        10'd612: TDATA = 37'b0100000001011111001000101100100001111;
        10'd613: TDATA = 37'b0100000000101101000011001100100000111;
        10'd614: TDATA = 37'b0011111111111011000001101100011111111;
        10'd615: TDATA = 37'b0011111111001001000100001100011111000;
        10'd616: TDATA = 37'b0011111110010111001010001100011110000;
        10'd617: TDATA = 37'b0011111101100101010100001100011101000;
        10'd618: TDATA = 37'b0011111100110011100010101100011100000;
        10'd619: TDATA = 37'b0011111100000001110100001100011011000;
        10'd620: TDATA = 37'b0011111011010000001010001100011010000;
        10'd621: TDATA = 37'b0011111010011110100011101100011001000;
        10'd622: TDATA = 37'b0011111001101101000001001100011000001;
        10'd623: TDATA = 37'b0011111000111011100010101100010111000;
        10'd624: TDATA = 37'b0011111000001010000111101100010110001;
        10'd625: TDATA = 37'b0011110111011000110000101100010101011;
        10'd626: TDATA = 37'b0011110110100111011101101100010100001;
        10'd627: TDATA = 37'b0011110101110110001110001100010011011;
        10'd628: TDATA = 37'b0011110101000101000010101100010010100;
        10'd629: TDATA = 37'b0011110100010011111011001100010001100;
        10'd630: TDATA = 37'b0011110011100010110111001100010000100;
        10'd631: TDATA = 37'b0011110010110001110110101100001111100;
        10'd632: TDATA = 37'b0011110010000000111010101100001110100;
        10'd633: TDATA = 37'b0011110001010000000010001100001101101;
        10'd634: TDATA = 37'b0011110000011111001101001100001100101;
        10'd635: TDATA = 37'b0011101111101110011100001100001011101;
        10'd636: TDATA = 37'b0011101110111101101110101100001010111;
        10'd637: TDATA = 37'b0011101110001101000101001100001010000;
        10'd638: TDATA = 37'b0011101101011100011111101100001001000;
        10'd639: TDATA = 37'b0011101100101011111101101100001000000;
        10'd640: TDATA = 37'b0011101011111011011111001100000111000;
        10'd641: TDATA = 37'b0011101011001011000100101100000110000;
        10'd642: TDATA = 37'b0011101010011010101101101100000101001;
        10'd643: TDATA = 37'b0011101001101010011010101100000100011;
        10'd644: TDATA = 37'b0011101000111010001011001100000011011;
        10'd645: TDATA = 37'b0011101000001001111111101100000010100;
        10'd646: TDATA = 37'b0011100111011001110111101100000001100;
        10'd647: TDATA = 37'b0011100110101001110011001100000000100;
        10'd648: TDATA = 37'b0011100101111001110010101011111111101;
        10'd649: TDATA = 37'b0011100101001001110101101011111110111;
        10'd650: TDATA = 37'b0011100100011001111100001011111101111;
        10'd651: TDATA = 37'b0011100011101010000110101011111101000;
        10'd652: TDATA = 37'b0011100010111010010100001011111100000;
        10'd653: TDATA = 37'b0011100010001010100110001011111011000;
        10'd654: TDATA = 37'b0011100001011010111011001011111010001;
        10'd655: TDATA = 37'b0011100000101011010100001011111001011;
        10'd656: TDATA = 37'b0011011111111011110000101011111000011;
        10'd657: TDATA = 37'b0011011111001100010000101011110111100;
        10'd658: TDATA = 37'b0011011110011100110100101011110110100;
        10'd659: TDATA = 37'b0011011101101101011100001011110101101;
        10'd660: TDATA = 37'b0011011100111110000110101011110100111;
        10'd661: TDATA = 37'b0011011100001110110101101011110011111;
        10'd662: TDATA = 37'b0011011011011111100111101011110011000;
        10'd663: TDATA = 37'b0011011010110000011101001011110010000;
        10'd664: TDATA = 37'b0011011010000001010110101011110001001;
        10'd665: TDATA = 37'b0011011001010010010011101011110000011;
        10'd666: TDATA = 37'b0011011000100011010011101011101111100;
        10'd667: TDATA = 37'b0011010111110100010111101011101110100;
        10'd668: TDATA = 37'b0011010111000101011111001011101101101;
        10'd669: TDATA = 37'b0011010110010110101010101011101100101;
        10'd670: TDATA = 37'b0011010101100111111001001011101011111;
        10'd671: TDATA = 37'b0011010100111001001011001011101011000;
        10'd672: TDATA = 37'b0011010100001010100000101011101010000;
        10'd673: TDATA = 37'b0011010011011011111010001011101001001;
        10'd674: TDATA = 37'b0011010010101101010110101011101000011;
        10'd675: TDATA = 37'b0011010001111110110111001011100111100;
        10'd676: TDATA = 37'b0011010001010000011010101011100110101;
        10'd677: TDATA = 37'b0011010000100010000001101011100101101;
        10'd678: TDATA = 37'b0011001111110011101100101011100100111;
        10'd679: TDATA = 37'b0011001111000101011010101011100100000;
        10'd680: TDATA = 37'b0011001110010111001100001011100011000;
        10'd681: TDATA = 37'b0011001101101001000001101011100010011;
        10'd682: TDATA = 37'b0011001100111010111010001011100001011;
        10'd683: TDATA = 37'b0011001100001100110110001011100000100;
        10'd684: TDATA = 37'b0011001011011110110101101011011111101;
        10'd685: TDATA = 37'b0011001010110000111000101011011110111;
        10'd686: TDATA = 37'b0011001010000010111110101011011110000;
        10'd687: TDATA = 37'b0011001001010101001000101011011101000;
        10'd688: TDATA = 37'b0011001000100111010101101011011100001;
        10'd689: TDATA = 37'b0011000111111001100110101011011011100;
        10'd690: TDATA = 37'b0011000111001011111010101011011010100;
        10'd691: TDATA = 37'b0011000110011110010010001011011001101;
        10'd692: TDATA = 37'b0011000101110000101101001011011000111;
        10'd693: TDATA = 37'b0011000101000011001011001011011000000;
        10'd694: TDATA = 37'b0011000100010101101100101011010111001;
        10'd695: TDATA = 37'b0011000011101000010001101011010110011;
        10'd696: TDATA = 37'b0011000010111010111010001011010101100;
        10'd697: TDATA = 37'b0011000010001101100110001011010100100;
        10'd698: TDATA = 37'b0011000001100000010101001011010011111;
        10'd699: TDATA = 37'b0011000000110011000111101011010011000;
        10'd700: TDATA = 37'b0011000000000101111101101011010010000;
        10'd701: TDATA = 37'b0010111111011000110111001011010001011;
        10'd702: TDATA = 37'b0010111110101011110011101011010000011;
        10'd703: TDATA = 37'b0010111101111110110011101011001111100;
        10'd704: TDATA = 37'b0010111101010001110110101011001110101;
        10'd705: TDATA = 37'b0010111100100100111101001011001110000;
        10'd706: TDATA = 37'b0010111011111000000111001011001101000;
        10'd707: TDATA = 37'b0010111011001011010100001011001100001;
        10'd708: TDATA = 37'b0010111010011110100100101011001011100;
        10'd709: TDATA = 37'b0010111001110001111000101011001010100;
        10'd710: TDATA = 37'b0010111001000101001111101011001001111;
        10'd711: TDATA = 37'b0010111000011000101010001011001001000;
        10'd712: TDATA = 37'b0010110111101100001000001011001000001;
        10'd713: TDATA = 37'b0010110110111111101000101011000111011;
        10'd714: TDATA = 37'b0010110110010011001101001011000110100;
        10'd715: TDATA = 37'b0010110101100110110100101011000101101;
        10'd716: TDATA = 37'b0010110100111010011111101011000100111;
        10'd717: TDATA = 37'b0010110100001110001101101011000100000;
        10'd718: TDATA = 37'b0010110011100001111110101011000011001;
        10'd719: TDATA = 37'b0010110010110101110011001011000010100;
        10'd720: TDATA = 37'b0010110010001001101011001011000001100;
        10'd721: TDATA = 37'b0010110001011101100110001011000000111;
        10'd722: TDATA = 37'b0010110000110001100100101011000000000;
        10'd723: TDATA = 37'b0010110000000101100110001010111111001;
        10'd724: TDATA = 37'b0010101111011001101010101010111110100;
        10'd725: TDATA = 37'b0010101110101101110010101010111101100;
        10'd726: TDATA = 37'b0010101110000001111101101010111100111;
        10'd727: TDATA = 37'b0010101101010110001100001010111100000;
        10'd728: TDATA = 37'b0010101100101010011101101010111011001;
        10'd729: TDATA = 37'b0010101011111110110010001010111010011;
        10'd730: TDATA = 37'b0010101011010011001010001010111001100;
        10'd731: TDATA = 37'b0010101010100111100101001010111000111;
        10'd732: TDATA = 37'b0010101001111100000011101010111000000;
        10'd733: TDATA = 37'b0010101001010000100101001010110111001;
        10'd734: TDATA = 37'b0010101000100101001001101010110110100;
        10'd735: TDATA = 37'b0010100111111001110001001010110101101;
        10'd736: TDATA = 37'b0010100111001110011100001010110100111;
        10'd737: TDATA = 37'b0010100110100011001010001010110100000;
        10'd738: TDATA = 37'b0010100101110111111011101010110011001;
        10'd739: TDATA = 37'b0010100101001100101111101010110010100;
        10'd740: TDATA = 37'b0010100100100001100111001010110001101;
        10'd741: TDATA = 37'b0010100011110110100001101010110001000;
        10'd742: TDATA = 37'b0010100011001011011111101010110000000;
        10'd743: TDATA = 37'b0010100010100000100000001010101111100;
        10'd744: TDATA = 37'b0010100001110101100100001010101110100;
        10'd745: TDATA = 37'b0010100001001010101011001010101101111;
        10'd746: TDATA = 37'b0010100000011111110101101010101101000;
        10'd747: TDATA = 37'b0010011111110101000010101010101100011;
        10'd748: TDATA = 37'b0010011111001010010011001010101011100;
        10'd749: TDATA = 37'b0010011110011111100110101010101010101;
        10'd750: TDATA = 37'b0010011101110100111101001010101010000;
        10'd751: TDATA = 37'b0010011101001010010110101010101001001;
        10'd752: TDATA = 37'b0010011100011111110011001010101000100;
        10'd753: TDATA = 37'b0010011011110101010011001010100111101;
        10'd754: TDATA = 37'b0010011011001010110101101010100110111;
        10'd755: TDATA = 37'b0010011010100000011011101010100110001;
        10'd756: TDATA = 37'b0010011001110110000100101010100101011;
        10'd757: TDATA = 37'b0010011001001011110000001010100100100;
        10'd758: TDATA = 37'b0010011000100001011111001010100011111;
        10'd759: TDATA = 37'b0010010111110111010001001010100011000;
        10'd760: TDATA = 37'b0010010111001101000110001010100010011;
        10'd761: TDATA = 37'b0010010110100010111110001010100001100;
        10'd762: TDATA = 37'b0010010101111000111001001010100000111;
        10'd763: TDATA = 37'b0010010101001110110111101010100000000;
        10'd764: TDATA = 37'b0010010100100100111000101010011111011;
        10'd765: TDATA = 37'b0010010011111010111100101010011110100;
        10'd766: TDATA = 37'b0010010011010001000011101010011101111;
        10'd767: TDATA = 37'b0010010010100111001101101010011101000;
        10'd768: TDATA = 37'b0010010001111101011010101010011100011;
        10'd769: TDATA = 37'b0010010001010011101010101010011011100;
        10'd770: TDATA = 37'b0010010000101001111110001010011010111;
        10'd771: TDATA = 37'b0010010000000000010100001010011010001;
        10'd772: TDATA = 37'b0010001111010110101100101010011001011;
        10'd773: TDATA = 37'b0010001110101101001000101010011000101;
        10'd774: TDATA = 37'b0010001110000011100111101010010111111;
        10'd775: TDATA = 37'b0010001101011010001001101010010111001;
        10'd776: TDATA = 37'b0010001100110000101110001010010110100;
        10'd777: TDATA = 37'b0010001100000111010110001010010101101;
        10'd778: TDATA = 37'b0010001011011110000000101010010101000;
        10'd779: TDATA = 37'b0010001010110100101110001010010100001;
        10'd780: TDATA = 37'b0010001010001011011110101010010011100;
        10'd781: TDATA = 37'b0010001001100010010010001010010010101;
        10'd782: TDATA = 37'b0010001000111001001000101010010010000;
        10'd783: TDATA = 37'b0010001000010000000010001010010001011;
        10'd784: TDATA = 37'b0010000111100110111110001010010000100;
        10'd785: TDATA = 37'b0010000110111101111101001010001111111;
        10'd786: TDATA = 37'b0010000110010100111111001010001111000;
        10'd787: TDATA = 37'b0010000101101100000100001010001110100;
        10'd788: TDATA = 37'b0010000101000011001100001010001101101;
        10'd789: TDATA = 37'b0010000100011010010110101010001101000;
        10'd790: TDATA = 37'b0010000011110001100100001010001100001;
        10'd791: TDATA = 37'b0010000011001000110100101010001011100;
        10'd792: TDATA = 37'b0010000010100000000111101010001010111;
        10'd793: TDATA = 37'b0010000001110111011110001010001010000;
        10'd794: TDATA = 37'b0010000001001110110111001010001001011;
        10'd795: TDATA = 37'b0010000000100110010011001010001000101;
        10'd796: TDATA = 37'b0001111111111101110001101010001000000;
        10'd797: TDATA = 37'b0001111111010101010011001010000111001;
        10'd798: TDATA = 37'b0001111110101100110111101010000110100;
        10'd799: TDATA = 37'b0001111110000100011111001010000101111;
        10'd800: TDATA = 37'b0001111101011100001001001010000101000;
        10'd801: TDATA = 37'b0001111100110011110110001010000100011;
        10'd802: TDATA = 37'b0001111100001011100101101010000011101;
        10'd803: TDATA = 37'b0001111011100011011000001010000011000;
        10'd804: TDATA = 37'b0001111010111011001101101010000010001;
        10'd805: TDATA = 37'b0001111010010011000101101010000001100;
        10'd806: TDATA = 37'b0001111001101011000000101010000000111;
        10'd807: TDATA = 37'b0001111001000010111110101010000000001;
        10'd808: TDATA = 37'b0001111000011010111111001001111111100;
        10'd809: TDATA = 37'b0001110111110011000010101001111110111;
        10'd810: TDATA = 37'b0001110111001011001000101001111110000;
        10'd811: TDATA = 37'b0001110110100011010001101001111101011;
        10'd812: TDATA = 37'b0001110101111011011101101001111100101;
        10'd813: TDATA = 37'b0001110101010011101100001001111100000;
        10'd814: TDATA = 37'b0001110100101011111101001001111011011;
        10'd815: TDATA = 37'b0001110100000100010001001001111010101;
        10'd816: TDATA = 37'b0001110011011100101000001001111010000;
        10'd817: TDATA = 37'b0001110010110101000001101001111001001;
        10'd818: TDATA = 37'b0001110010001101011110001001111000100;
        10'd819: TDATA = 37'b0001110001100101111101001001110111111;
        10'd820: TDATA = 37'b0001110000111110011110101001110111001;
        10'd821: TDATA = 37'b0001110000010111000011001001110110100;
        10'd822: TDATA = 37'b0001101111101111101010101001110101111;
        10'd823: TDATA = 37'b0001101111001000010100101001110101001;
        10'd824: TDATA = 37'b0001101110100001000001001001110100100;
        10'd825: TDATA = 37'b0001101101111001110000101001110011111;
        10'd826: TDATA = 37'b0001101101010010100011001001110011000;
        10'd827: TDATA = 37'b0001101100101011010111101001110010100;
        10'd828: TDATA = 37'b0001101100000100001111101001110001111;
        10'd829: TDATA = 37'b0001101011011101001001101001110001000;
        10'd830: TDATA = 37'b0001101010110110000110101001110000100;
        10'd831: TDATA = 37'b0001101010001111000110001001101111101;
        10'd832: TDATA = 37'b0001101001101000001000101001101111000;
        10'd833: TDATA = 37'b0001101001000001001101101001101110100;
        10'd834: TDATA = 37'b0001101000011010010101101001101101101;
        10'd835: TDATA = 37'b0001100111110011011111101001101101000;
        10'd836: TDATA = 37'b0001100111001100101101001001101100100;
        10'd837: TDATA = 37'b0001100110100101111100101001101011101;
        10'd838: TDATA = 37'b0001100101111111001111001001101011000;
        10'd839: TDATA = 37'b0001100101011000100100001001101010100;
        10'd840: TDATA = 37'b0001100100110001111011101001101001101;
        10'd841: TDATA = 37'b0001100100001011010110001001101001000;
        10'd842: TDATA = 37'b0001100011100100110011001001101000100;
        10'd843: TDATA = 37'b0001100010111110010010101001100111101;
        10'd844: TDATA = 37'b0001100010010111110101001001100111000;
        10'd845: TDATA = 37'b0001100001110001011010001001100110100;
        10'd846: TDATA = 37'b0001100001001011000001101001100101101;
        10'd847: TDATA = 37'b0001100000100100101011101001100101000;
        10'd848: TDATA = 37'b0001011111111110011000101001100100100;
        10'd849: TDATA = 37'b0001011111011000001000001001100011111;
        10'd850: TDATA = 37'b0001011110110001111010001001100011001;
        10'd851: TDATA = 37'b0001011110001011101110101001100010100;
        10'd852: TDATA = 37'b0001011101100101100110001001100001111;
        10'd853: TDATA = 37'b0001011100111111011111101001100001001;
        10'd854: TDATA = 37'b0001011100011001011100001001100000100;
        10'd855: TDATA = 37'b0001011011110011011011001001011111111;
        10'd856: TDATA = 37'b0001011011001101011101001001011111001;
        10'd857: TDATA = 37'b0001011010100111100001001001011110100;
        10'd858: TDATA = 37'b0001011010000001101000001001011110000;
        10'd859: TDATA = 37'b0001011001011011110001001001011101011;
        10'd860: TDATA = 37'b0001011000110101111101001001011100101;
        10'd861: TDATA = 37'b0001011000010000001011101001011100000;
        10'd862: TDATA = 37'b0001010111101010011100101001011011011;
        10'd863: TDATA = 37'b0001010111000100110000001001011010111;
        10'd864: TDATA = 37'b0001010110011111000110101001011010000;
        10'd865: TDATA = 37'b0001010101111001011111001001011001100;
        10'd866: TDATA = 37'b0001010101010011111010101001011000111;
        10'd867: TDATA = 37'b0001010100101110011000001001011000001;
        10'd868: TDATA = 37'b0001010100001000111000101001010111100;
        10'd869: TDATA = 37'b0001010011100011011011101001010111000;
        10'd870: TDATA = 37'b0001010010111110000001001001010110011;
        10'd871: TDATA = 37'b0001010010011000101001001001010101101;
        10'd872: TDATA = 37'b0001010001110011010011101001010101000;
        10'd873: TDATA = 37'b0001010001001110000000101001010100100;
        10'd874: TDATA = 37'b0001010000101000110000001001010011111;
        10'd875: TDATA = 37'b0001010000000011100010001001010011001;
        10'd876: TDATA = 37'b0001001111011110010110101001010010100;
        10'd877: TDATA = 37'b0001001110111001001101101001010010000;
        10'd878: TDATA = 37'b0001001110010100000111001001010001011;
        10'd879: TDATA = 37'b0001001101101111000011001001010000101;
        10'd880: TDATA = 37'b0001001101001010000001101001010000000;
        10'd881: TDATA = 37'b0001001100100101000010101001001111100;
        10'd882: TDATA = 37'b0001001100000000000110001001001110111;
        10'd883: TDATA = 37'b0001001011011011001100001001001110001;
        10'd884: TDATA = 37'b0001001010110110010100001001001101100;
        10'd885: TDATA = 37'b0001001010010001011111001001001101000;
        10'd886: TDATA = 37'b0001001001101100101100101001001100011;
        10'd887: TDATA = 37'b0001001001000111111100101001001011101;
        10'd888: TDATA = 37'b0001001000100011001110101001001011000;
        10'd889: TDATA = 37'b0001000111111110100011101001001010100;
        10'd890: TDATA = 37'b0001000111011001111010101001001001111;
        10'd891: TDATA = 37'b0001000110110101010100001001001001011;
        10'd892: TDATA = 37'b0001000110010000110000101001001000101;
        10'd893: TDATA = 37'b0001000101101100001111001001001000000;
        10'd894: TDATA = 37'b0001000101000111110000001001000111100;
        10'd895: TDATA = 37'b0001000100100011010011001001000110111;
        10'd896: TDATA = 37'b0001000011111110111001001001000110001;
        10'd897: TDATA = 37'b0001000011011010100001001001000101100;
        10'd898: TDATA = 37'b0001000010110110001100001001000101000;
        10'd899: TDATA = 37'b0001000010010001111001001001000100100;
        10'd900: TDATA = 37'b0001000001101101101000101001000011111;
        10'd901: TDATA = 37'b0001000001001001011010101001000011001;
        10'd902: TDATA = 37'b0001000000100101001111001001000010100;
        10'd903: TDATA = 37'b0001000000000001000101101001000010000;
        10'd904: TDATA = 37'b0000111111011100111110101001000001100;
        10'd905: TDATA = 37'b0000111110111000111010001001000000111;
        10'd906: TDATA = 37'b0000111110010100111000001001000000001;
        10'd907: TDATA = 37'b0000111101110000111000101000111111100;
        10'd908: TDATA = 37'b0000111101001100111011001000111111000;
        10'd909: TDATA = 37'b0000111100101001000000001000111110100;
        10'd910: TDATA = 37'b0000111100000101000111101000111101111;
        10'd911: TDATA = 37'b0000111011100001010001101000111101001;
        10'd912: TDATA = 37'b0000111010111101011101101000111100101;
        10'd913: TDATA = 37'b0000111010011001101100001000111100000;
        10'd914: TDATA = 37'b0000111001110101111101001000111011100;
        10'd915: TDATA = 37'b0000111001010010010000101000111010111;
        10'd916: TDATA = 37'b0000111000101110100110001000111010011;
        10'd917: TDATA = 37'b0000111000001010111110001000111001101;
        10'd918: TDATA = 37'b0000110111100111011000101000111001000;
        10'd919: TDATA = 37'b0000110111000011110101001000111000100;
        10'd920: TDATA = 37'b0000110110100000010100001000111000000;
        10'd921: TDATA = 37'b0000110101111100110101101000110111011;
        10'd922: TDATA = 37'b0000110101011001011001001000110110111;
        10'd923: TDATA = 37'b0000110100110101111111001000110110001;
        10'd924: TDATA = 37'b0000110100010010100111101000110101100;
        10'd925: TDATA = 37'b0000110011101111010010001000110101000;
        10'd926: TDATA = 37'b0000110011001011111111001000110100100;
        10'd927: TDATA = 37'b0000110010101000101110001000110100000;
        10'd928: TDATA = 37'b0000110010000101100000001000110011011;
        10'd929: TDATA = 37'b0000110001100010010011101000110010101;
        10'd930: TDATA = 37'b0000110000111111001010001000110010000;
        10'd931: TDATA = 37'b0000110000011100000010101000110001100;
        10'd932: TDATA = 37'b0000101111111000111101101000110001000;
        10'd933: TDATA = 37'b0000101111010101111010101000110000100;
        10'd934: TDATA = 37'b0000101110110010111010001000101111111;
        10'd935: TDATA = 37'b0000101110001111111011101000101111001;
        10'd936: TDATA = 37'b0000101101101100111111101000101110101;
        10'd937: TDATA = 37'b0000101101001010000101101000101110000;
        10'd938: TDATA = 37'b0000101100100111001110001000101101100;
        10'd939: TDATA = 37'b0000101100000100011001001000101101000;
        10'd940: TDATA = 37'b0000101011100001100110001000101100100;
        10'd941: TDATA = 37'b0000101010111110110101101000101011111;
        10'd942: TDATA = 37'b0000101010011100000111001000101011011;
        10'd943: TDATA = 37'b0000101001111001011011001000101010101;
        10'd944: TDATA = 37'b0000101001010110110001001000101010001;
        10'd945: TDATA = 37'b0000101000110100001001101000101001101;
        10'd946: TDATA = 37'b0000101000010001100100001000101001000;
        10'd947: TDATA = 37'b0000100111101111000001001000101000100;
        10'd948: TDATA = 37'b0000100111001100100000001000101000000;
        10'd949: TDATA = 37'b0000100110101010000001101000100111011;
        10'd950: TDATA = 37'b0000100110000111100101001000100110111;
        10'd951: TDATA = 37'b0000100101100101001010101000100110011;
        10'd952: TDATA = 37'b0000100101000010110010101000100101101;
        10'd953: TDATA = 37'b0000100100100000011101001000100101001;
        10'd954: TDATA = 37'b0000100011111110001001101000100100100;
        10'd955: TDATA = 37'b0000100011011011111000001000100100000;
        10'd956: TDATA = 37'b0000100010111001101001001000100011100;
        10'd957: TDATA = 37'b0000100010010111011100001000100011000;
        10'd958: TDATA = 37'b0000100001110101010001101000100010011;
        10'd959: TDATA = 37'b0000100001010011001001001000100001111;
        10'd960: TDATA = 37'b0000100000110001000011001000100001011;
        10'd961: TDATA = 37'b0000100000001110111110101000100000101;
        10'd962: TDATA = 37'b0000011111101100111101001000100000001;
        10'd963: TDATA = 37'b0000011111001010111101001000011111100;
        10'd964: TDATA = 37'b0000011110101000111111101000011111000;
        10'd965: TDATA = 37'b0000011110000111000100101000011110100;
        10'd966: TDATA = 37'b0000011101100101001011101000011110000;
        10'd967: TDATA = 37'b0000011101000011010100101000011101100;
        10'd968: TDATA = 37'b0000011100100001011111101000011101000;
        10'd969: TDATA = 37'b0000011011111111101101001000011100011;
        10'd970: TDATA = 37'b0000011011011101111100101000011011111;
        10'd971: TDATA = 37'b0000011010111100001110101000011011011;
        10'd972: TDATA = 37'b0000011010011010100010001000011010101;
        10'd973: TDATA = 37'b0000011001111000111000001000011010001;
        10'd974: TDATA = 37'b0000011001010111010000101000011001101;
        10'd975: TDATA = 37'b0000011000110101101011001000011001000;
        10'd976: TDATA = 37'b0000011000010100000111101000011000100;
        10'd977: TDATA = 37'b0000010111110010100110001000011000000;
        10'd978: TDATA = 37'b0000010111010001000111001000010111100;
        10'd979: TDATA = 37'b0000010110101111101001101000010111000;
        10'd980: TDATA = 37'b0000010110001110001111001000010110100;
        10'd981: TDATA = 37'b0000010101101100110110001000010110000;
        10'd982: TDATA = 37'b0000010101001011011111101000010101011;
        10'd983: TDATA = 37'b0000010100101010001011001000010100111;
        10'd984: TDATA = 37'b0000010100001000111000101000010100011;
        10'd985: TDATA = 37'b0000010011100111101000001000010011101;
        10'd986: TDATA = 37'b0000010011000110011010001000010011001;
        10'd987: TDATA = 37'b0000010010100101001110001000010010101;
        10'd988: TDATA = 37'b0000010010000100000100001000010010001;
        10'd989: TDATA = 37'b0000010001100010111100001000010001101;
        10'd990: TDATA = 37'b0000010001000001110110101000010001001;
        10'd991: TDATA = 37'b0000010000100000110011001000010000101;
        10'd992: TDATA = 37'b0000001111111111110001101000010000000;
        10'd993: TDATA = 37'b0000001111011110110010001000001111100;
        10'd994: TDATA = 37'b0000001110111101110100101000001111000;
        10'd995: TDATA = 37'b0000001110011100111001001000001110100;
        10'd996: TDATA = 37'b0000001101111100000000001000001110000;
        10'd997: TDATA = 37'b0000001101011011001001001000001101100;
        10'd998: TDATA = 37'b0000001100111010010100001000001101000;
        10'd999: TDATA = 37'b0000001100011001100001001000001100100;
        10'd1000: TDATA = 37'b0000001011111000110000001000001100000;
        10'd1001: TDATA = 37'b0000001011011000000001101000001011100;
        10'd1002: TDATA = 37'b0000001010110111010100101000001010111;
        10'd1003: TDATA = 37'b0000001010010110101010001000001010011;
        10'd1004: TDATA = 37'b0000001001110110000001101000001001111;
        10'd1005: TDATA = 37'b0000001001010101011011001000001001011;
        10'd1006: TDATA = 37'b0000001000110100110110101000001000111;
        10'd1007: TDATA = 37'b0000001000010100010100001000001000011;
        10'd1008: TDATA = 37'b0000000111110011110011101000000111111;
        10'd1009: TDATA = 37'b0000000111010011010101001000000111011;
        10'd1010: TDATA = 37'b0000000110110010111001001000000110111;
        10'd1011: TDATA = 37'b0000000110010010011110101000000110011;
        10'd1012: TDATA = 37'b0000000101110010000110101000000101111;
        10'd1013: TDATA = 37'b0000000101010001110000101000000101011;
        10'd1014: TDATA = 37'b0000000100110001011100001000000100111;
        10'd1015: TDATA = 37'b0000000100010001001010001000000100011;
        10'd1016: TDATA = 37'b0000000011110000111010001000000011111;
        10'd1017: TDATA = 37'b0000000011010000101100001000000011011;
        10'd1018: TDATA = 37'b0000000010110000100000001000000010111;
        10'd1019: TDATA = 37'b0000000010010000010110001000000010011;
        10'd1020: TDATA = 37'b0000000001110000001110001000000001111;
        10'd1021: TDATA = 37'b0000000001010000001000001000000001011;
        10'd1022: TDATA = 37'b0000000000110000000100001000000000111;
        10'd1023: TDATA = 37'b0000000000010000000010001000000000011;
        endcase
    end
    endfunction

    wire sx;
    wire [7:0] ex;
    assign sx = x[31];
    assign ex = x[30:23];

    // pm = 1 のとき - 0のとき +
    wire [9:0] ml;
    wire pm;
    wire [11:0] mr;
    assign ml = x[22:13];
    assign pm = x[12];
    assign mr = x[11:0];

    wire [36:0] tdata;
    assign tdata = TDATA(ml);

    wire [22:0] a0_inv;
    wire [13:0] a02_inv;
    assign a0_inv = tdata[36:14];
    assign a02_inv = tdata[13:0];

    wire [11:0] notmr;
    assign notmr = ~mr;

    wire [35:0] my_extend1;
    assign my_extend1 = {a0_inv,13'b0} - mr * a02_inv;

    wire [35:0] my_extend2;
    assign my_extend2 = {a0_inv,13'b0} + notmr * a02_inv;

    wire [22:0] my;
    assign my = (pm) ? my_extend1[35:13]: my_extend2[35:13];

    wire [8:0] eya;
    assign eya = 9'd253 - ex;

    wire [7:0] ey;
    assign ey = (eya[8]) ? 0: eya[7:0];

    assign y = {sx,ey,my};

endmodule

