module fsqrt(
    input wire [31:0] x,
    output wire [31:0] y);

    function [36:0] TDATA (
	input [10:0] KEY
    );
    begin
        case(KEY)
        11'd1024: TDATA = 37'b0000000000000000000000010000000000000;
        11'd1025: TDATA = 37'b0000000000011111111111101111111111100;
        11'd1026: TDATA = 37'b0000000000111111111110001111111111000;
        11'd1027: TDATA = 37'b0000000001011111111011101111111110100;
        11'd1028: TDATA = 37'b0000000001111111111000001111111110000;
        11'd1029: TDATA = 37'b0000000010011111110011101111111101100;
        11'd1030: TDATA = 37'b0000000010111111101110001111111101000;
        11'd1031: TDATA = 37'b0000000011011111100111101111111100100;
        11'd1032: TDATA = 37'b0000000011111111100000001111111100000;
        11'd1033: TDATA = 37'b0000000100011111010111101111111011100;
        11'd1034: TDATA = 37'b0000000100111111001110001111111011000;
        11'd1035: TDATA = 37'b0000000101011111000100001111111010100;
        11'd1036: TDATA = 37'b0000000101111110111000101111111010000;
        11'd1037: TDATA = 37'b0000000110011110101100001111111001100;
        11'd1038: TDATA = 37'b0000000110111110011110101111111001001;
        11'd1039: TDATA = 37'b0000000111011110010000101111111000101;
        11'd1040: TDATA = 37'b0000000111111110000001001111111000001;
        11'd1041: TDATA = 37'b0000001000011101110000101111110111101;
        11'd1042: TDATA = 37'b0000001000111101011111101111110111001;
        11'd1043: TDATA = 37'b0000001001011101001101001111110110101;
        11'd1044: TDATA = 37'b0000001001111100111010001111110110001;
        11'd1045: TDATA = 37'b0000001010011100100101101111110101101;
        11'd1046: TDATA = 37'b0000001010111100010000101111110101001;
        11'd1047: TDATA = 37'b0000001011011011111010101111110100110;
        11'd1048: TDATA = 37'b0000001011111011100011101111110100010;
        11'd1049: TDATA = 37'b0000001100011011001011101111110011110;
        11'd1050: TDATA = 37'b0000001100111010110010001111110011010;
        11'd1051: TDATA = 37'b0000001101011010011000001111110010110;
        11'd1052: TDATA = 37'b0000001101111001111101101111110010010;
        11'd1053: TDATA = 37'b0000001110011001100001101111110001110;
        11'd1054: TDATA = 37'b0000001110111001000100101111110001011;
        11'd1055: TDATA = 37'b0000001111011000100110101111110000111;
        11'd1056: TDATA = 37'b0000001111111000001000001111110000011;
        11'd1057: TDATA = 37'b0000010000010111101000001111101111111;
        11'd1058: TDATA = 37'b0000010000110111000111101111101111011;
        11'd1059: TDATA = 37'b0000010001010110100101101111101110111;
        11'd1060: TDATA = 37'b0000010001110110000011001111101110100;
        11'd1061: TDATA = 37'b0000010010010101011111101111101110000;
        11'd1062: TDATA = 37'b0000010010110100111011001111101101100;
        11'd1063: TDATA = 37'b0000010011010100010101101111101101000;
        11'd1064: TDATA = 37'b0000010011110011101111101111101100101;
        11'd1065: TDATA = 37'b0000010100010011001000001111101100001;
        11'd1066: TDATA = 37'b0000010100110010011111101111101011101;
        11'd1067: TDATA = 37'b0000010101010001110110101111101011001;
        11'd1068: TDATA = 37'b0000010101110001001100101111101010101;
        11'd1069: TDATA = 37'b0000010110010000100001001111101010010;
        11'd1070: TDATA = 37'b0000010110101111110101001111101001110;
        11'd1071: TDATA = 37'b0000010111001111001000001111101001010;
        11'd1072: TDATA = 37'b0000010111101110011010001111101000110;
        11'd1073: TDATA = 37'b0000011000001101101011101111101000011;
        11'd1074: TDATA = 37'b0000011000101100111011101111100111111;
        11'd1075: TDATA = 37'b0000011001001100001011001111100111011;
        11'd1076: TDATA = 37'b0000011001101011011001101111100111000;
        11'd1077: TDATA = 37'b0000011010001010100110101111100110100;
        11'd1078: TDATA = 37'b0000011010101001110011001111100110000;
        11'd1079: TDATA = 37'b0000011011001000111111001111100101100;
        11'd1080: TDATA = 37'b0000011011101000001001101111100101001;
        11'd1081: TDATA = 37'b0000011100000111010011001111100100101;
        11'd1082: TDATA = 37'b0000011100100110011100001111100100001;
        11'd1083: TDATA = 37'b0000011101000101100100001111100011110;
        11'd1084: TDATA = 37'b0000011101100100101011001111100011010;
        11'd1085: TDATA = 37'b0000011110000011110001001111100010110;
        11'd1086: TDATA = 37'b0000011110100010110110001111100010011;
        11'd1087: TDATA = 37'b0000011111000001111010101111100001111;
        11'd1088: TDATA = 37'b0000011111100000111101101111100001011;
        11'd1089: TDATA = 37'b0000100000000000000000001111100001000;
        11'd1090: TDATA = 37'b0000100000011111000001101111100000100;
        11'd1091: TDATA = 37'b0000100000111110000010001111100000000;
        11'd1092: TDATA = 37'b0000100001011101000001101111011111101;
        11'd1093: TDATA = 37'b0000100001111100000000101111011111001;
        11'd1094: TDATA = 37'b0000100010011010111110101111011110110;
        11'd1095: TDATA = 37'b0000100010111001111011101111011110010;
        11'd1096: TDATA = 37'b0000100011011000110111101111011101110;
        11'd1097: TDATA = 37'b0000100011110111110010101111011101011;
        11'd1098: TDATA = 37'b0000100100010110101100101111011100111;
        11'd1099: TDATA = 37'b0000100100110101100110001111011100100;
        11'd1100: TDATA = 37'b0000100101010100011110101111011100000;
        11'd1101: TDATA = 37'b0000100101110011010110001111011011100;
        11'd1102: TDATA = 37'b0000100110010010001100101111011011001;
        11'd1103: TDATA = 37'b0000100110110001000010101111011010101;
        11'd1104: TDATA = 37'b0000100111001111110111001111011010010;
        11'd1105: TDATA = 37'b0000100111101110101011001111011001110;
        11'd1106: TDATA = 37'b0000101000001101011110001111011001010;
        11'd1107: TDATA = 37'b0000101000101100010000101111011000111;
        11'd1108: TDATA = 37'b0000101001001011000001101111011000011;
        11'd1109: TDATA = 37'b0000101001101001110010001111011000000;
        11'd1110: TDATA = 37'b0000101010001000100001101111010111100;
        11'd1111: TDATA = 37'b0000101010100111010000001111010111001;
        11'd1112: TDATA = 37'b0000101011000101111110001111010110101;
        11'd1113: TDATA = 37'b0000101011100100101011001111010110010;
        11'd1114: TDATA = 37'b0000101100000011010111001111010101110;
        11'd1115: TDATA = 37'b0000101100100010000010001111010101011;
        11'd1116: TDATA = 37'b0000101101000000101100001111010100111;
        11'd1117: TDATA = 37'b0000101101011111010101101111010100100;
        11'd1118: TDATA = 37'b0000101101111101111110001111010100000;
        11'd1119: TDATA = 37'b0000101110011100100101101111010011101;
        11'd1120: TDATA = 37'b0000101110111011001100001111010011001;
        11'd1121: TDATA = 37'b0000101111011001110010001111010010110;
        11'd1122: TDATA = 37'b0000101111111000010111001111010010010;
        11'd1123: TDATA = 37'b0000110000010110111011001111010001111;
        11'd1124: TDATA = 37'b0000110000110101011110001111010001011;
        11'd1125: TDATA = 37'b0000110001010100000000101111010001000;
        11'd1126: TDATA = 37'b0000110001110010100010001111010000100;
        11'd1127: TDATA = 37'b0000110010010001000010101111010000001;
        11'd1128: TDATA = 37'b0000110010101111100010101111001111101;
        11'd1129: TDATA = 37'b0000110011001110000001001111001111010;
        11'd1130: TDATA = 37'b0000110011101100011111001111001110110;
        11'd1131: TDATA = 37'b0000110100001010111100101111001110011;
        11'd1132: TDATA = 37'b0000110100101001011000101111001101111;
        11'd1133: TDATA = 37'b0000110101000111110100001111001101100;
        11'd1134: TDATA = 37'b0000110101100110001110101111001101001;
        11'd1135: TDATA = 37'b0000110110000100101000101111001100101;
        11'd1136: TDATA = 37'b0000110110100011000001001111001100010;
        11'd1137: TDATA = 37'b0000110111000001011001001111001011110;
        11'd1138: TDATA = 37'b0000110111011111110000101111001011011;
        11'd1139: TDATA = 37'b0000110111111110000110101111001010111;
        11'd1140: TDATA = 37'b0000111000011100011100001111001010100;
        11'd1141: TDATA = 37'b0000111000111010110000101111001010001;
        11'd1142: TDATA = 37'b0000111001011001000100101111001001101;
        11'd1143: TDATA = 37'b0000111001110111010111101111001001010;
        11'd1144: TDATA = 37'b0000111010010101101001101111001000110;
        11'd1145: TDATA = 37'b0000111010110011111010101111001000011;
        11'd1146: TDATA = 37'b0000111011010010001011001111001000000;
        11'd1147: TDATA = 37'b0000111011110000011010101111000111100;
        11'd1148: TDATA = 37'b0000111100001110101001001111000111001;
        11'd1149: TDATA = 37'b0000111100101100110111001111000110110;
        11'd1150: TDATA = 37'b0000111101001011000100001111000110010;
        11'd1151: TDATA = 37'b0000111101101001010000001111000101111;
        11'd1152: TDATA = 37'b0000111110000111011011001111000101011;
        11'd1153: TDATA = 37'b0000111110100101100101101111000101000;
        11'd1154: TDATA = 37'b0000111111000011101111101111000100101;
        11'd1155: TDATA = 37'b0000111111100001111000001111000100001;
        11'd1156: TDATA = 37'b0001000000000000000000001111000011110;
        11'd1157: TDATA = 37'b0001000000011110000111001111000011011;
        11'd1158: TDATA = 37'b0001000000111100001101101111000010111;
        11'd1159: TDATA = 37'b0001000001011010010011001111000010100;
        11'd1160: TDATA = 37'b0001000001111000010111101111000010001;
        11'd1161: TDATA = 37'b0001000010010110011011001111000001101;
        11'd1162: TDATA = 37'b0001000010110100011110001111000001010;
        11'd1163: TDATA = 37'b0001000011010010100000101111000000111;
        11'd1164: TDATA = 37'b0001000011110000100001101111000000100;
        11'd1165: TDATA = 37'b0001000100001110100010001111000000000;
        11'd1166: TDATA = 37'b0001000100101100100010001110111111101;
        11'd1167: TDATA = 37'b0001000101001010100000101110111111010;
        11'd1168: TDATA = 37'b0001000101101000011110101110111110110;
        11'd1169: TDATA = 37'b0001000110000110011100001110111110011;
        11'd1170: TDATA = 37'b0001000110100100011000001110111110000;
        11'd1171: TDATA = 37'b0001000111000010010100001110111101101;
        11'd1172: TDATA = 37'b0001000111100000001110101110111101001;
        11'd1173: TDATA = 37'b0001000111111110001000101110111100110;
        11'd1174: TDATA = 37'b0001001000011100000001101110111100011;
        11'd1175: TDATA = 37'b0001001000111001111010001110111100000;
        11'd1176: TDATA = 37'b0001001001010111110001101110111011100;
        11'd1177: TDATA = 37'b0001001001110101101000001110111011001;
        11'd1178: TDATA = 37'b0001001010010011011110001110111010110;
        11'd1179: TDATA = 37'b0001001010110001010011001110111010011;
        11'd1180: TDATA = 37'b0001001011001111000111001110111001111;
        11'd1181: TDATA = 37'b0001001011101100111010101110111001100;
        11'd1182: TDATA = 37'b0001001100001010101101001110111001001;
        11'd1183: TDATA = 37'b0001001100101000011111001110111000110;
        11'd1184: TDATA = 37'b0001001101000110010000001110111000010;
        11'd1185: TDATA = 37'b0001001101100100000000001110110111111;
        11'd1186: TDATA = 37'b0001001110000001101111101110110111100;
        11'd1187: TDATA = 37'b0001001110011111011110001110110111001;
        11'd1188: TDATA = 37'b0001001110111101001100001110110110110;
        11'd1189: TDATA = 37'b0001001111011010111001001110110110010;
        11'd1190: TDATA = 37'b0001001111111000100101001110110101111;
        11'd1191: TDATA = 37'b0001010000010110010000101110110101100;
        11'd1192: TDATA = 37'b0001010000110011111011001110110101001;
        11'd1193: TDATA = 37'b0001010001010001100101001110110100110;
        11'd1194: TDATA = 37'b0001010001101111001110001110110100010;
        11'd1195: TDATA = 37'b0001010010001100110110001110110011111;
        11'd1196: TDATA = 37'b0001010010101010011101101110110011100;
        11'd1197: TDATA = 37'b0001010011001000000100001110110011001;
        11'd1198: TDATA = 37'b0001010011100101101010001110110010110;
        11'd1199: TDATA = 37'b0001010100000011001111001110110010011;
        11'd1200: TDATA = 37'b0001010100100000110011101110110001111;
        11'd1201: TDATA = 37'b0001010100111110010110101110110001100;
        11'd1202: TDATA = 37'b0001010101011011111001101110110001001;
        11'd1203: TDATA = 37'b0001010101111001011011101110110000110;
        11'd1204: TDATA = 37'b0001010110010110111100101110110000011;
        11'd1205: TDATA = 37'b0001010110110100011100101110110000000;
        11'd1206: TDATA = 37'b0001010111010001111100101110101111101;
        11'd1207: TDATA = 37'b0001010111101111011011001110101111001;
        11'd1208: TDATA = 37'b0001011000001100111001001110101110110;
        11'd1209: TDATA = 37'b0001011000101010010110001110101110011;
        11'd1210: TDATA = 37'b0001011001000111110010101110101110000;
        11'd1211: TDATA = 37'b0001011001100101001110101110101101101;
        11'd1212: TDATA = 37'b0001011010000010101001001110101101010;
        11'd1213: TDATA = 37'b0001011010100000000011001110101100111;
        11'd1214: TDATA = 37'b0001011010111101011100101110101100100;
        11'd1215: TDATA = 37'b0001011011011010110101001110101100001;
        11'd1216: TDATA = 37'b0001011011111000001101001110101011101;
        11'd1217: TDATA = 37'b0001011100010101100100001110101011010;
        11'd1218: TDATA = 37'b0001011100110010111010001110101010111;
        11'd1219: TDATA = 37'b0001011101010000001111101110101010100;
        11'd1220: TDATA = 37'b0001011101101101100100001110101010001;
        11'd1221: TDATA = 37'b0001011110001010111000001110101001110;
        11'd1222: TDATA = 37'b0001011110101000001011001110101001011;
        11'd1223: TDATA = 37'b0001011111000101011101101110101001000;
        11'd1224: TDATA = 37'b0001011111100010101111001110101000101;
        11'd1225: TDATA = 37'b0001100000000000000000001110101000010;
        11'd1226: TDATA = 37'b0001100000011101010000001110100111111;
        11'd1227: TDATA = 37'b0001100000111010011111101110100111100;
        11'd1228: TDATA = 37'b0001100001010111101110001110100111001;
        11'd1229: TDATA = 37'b0001100001110100111011101110100110110;
        11'd1230: TDATA = 37'b0001100010010010001001001110100110011;
        11'd1231: TDATA = 37'b0001100010101111010101001110100110000;
        11'd1232: TDATA = 37'b0001100011001100100000101110100101101;
        11'd1233: TDATA = 37'b0001100011101001101011101110100101001;
        11'd1234: TDATA = 37'b0001100100000110110101101110100100110;
        11'd1235: TDATA = 37'b0001100100100011111110101110100100011;
        11'd1236: TDATA = 37'b0001100101000001000111001110100100000;
        11'd1237: TDATA = 37'b0001100101011110001110101110100011101;
        11'd1238: TDATA = 37'b0001100101111011010101101110100011010;
        11'd1239: TDATA = 37'b0001100110011000011100001110100010111;
        11'd1240: TDATA = 37'b0001100110110101100001101110100010100;
        11'd1241: TDATA = 37'b0001100111010010100110001110100010001;
        11'd1242: TDATA = 37'b0001100111101111101010001110100001110;
        11'd1243: TDATA = 37'b0001101000001100101101101110100001011;
        11'd1244: TDATA = 37'b0001101000101001110000001110100001000;
        11'd1245: TDATA = 37'b0001101001000110110001101110100000101;
        11'd1246: TDATA = 37'b0001101001100011110010101110100000010;
        11'd1247: TDATA = 37'b0001101010000000110010101110011111111;
        11'd1248: TDATA = 37'b0001101010011101110010001110011111100;
        11'd1249: TDATA = 37'b0001101010111010110001001110011111010;
        11'd1250: TDATA = 37'b0001101011010111101111001110011110111;
        11'd1251: TDATA = 37'b0001101011110100101100101110011110100;
        11'd1252: TDATA = 37'b0001101100010001101001001110011110001;
        11'd1253: TDATA = 37'b0001101100101110100100101110011101110;
        11'd1254: TDATA = 37'b0001101101001011011111101110011101011;
        11'd1255: TDATA = 37'b0001101101101000011010001110011101000;
        11'd1256: TDATA = 37'b0001101110000101010011101110011100101;
        11'd1257: TDATA = 37'b0001101110100010001100101110011100010;
        11'd1258: TDATA = 37'b0001101110111111000100101110011011111;
        11'd1259: TDATA = 37'b0001101111011011111100001110011011100;
        11'd1260: TDATA = 37'b0001101111111000110010101110011011001;
        11'd1261: TDATA = 37'b0001110000010101101000101110011010110;
        11'd1262: TDATA = 37'b0001110000110010011101101110011010011;
        11'd1263: TDATA = 37'b0001110001001111010010001110011010000;
        11'd1264: TDATA = 37'b0001110001101100000101101110011001101;
        11'd1265: TDATA = 37'b0001110010001000111000101110011001010;
        11'd1266: TDATA = 37'b0001110010100101101011001110011001000;
        11'd1267: TDATA = 37'b0001110011000010011100101110011000101;
        11'd1268: TDATA = 37'b0001110011011111001101001110011000010;
        11'd1269: TDATA = 37'b0001110011111011111101101110010111111;
        11'd1270: TDATA = 37'b0001110100011000101100101110010111100;
        11'd1271: TDATA = 37'b0001110100110101011011101110010111001;
        11'd1272: TDATA = 37'b0001110101010010001001001110010110110;
        11'd1273: TDATA = 37'b0001110101101110110110101110010110011;
        11'd1274: TDATA = 37'b0001110110001011100011001110010110000;
        11'd1275: TDATA = 37'b0001110110101000001110101110010101110;
        11'd1276: TDATA = 37'b0001110111000100111001101110010101011;
        11'd1277: TDATA = 37'b0001110111100001100100001110010101000;
        11'd1278: TDATA = 37'b0001110111111110001101101110010100101;
        11'd1279: TDATA = 37'b0001111000011010110110101110010100010;
        11'd1280: TDATA = 37'b0001111000110111011110101110010011111;
        11'd1281: TDATA = 37'b0001111001010100000110001110010011100;
        11'd1282: TDATA = 37'b0001111001110000101100101110010011001;
        11'd1283: TDATA = 37'b0001111010001101010010101110010010111;
        11'd1284: TDATA = 37'b0001111010101001111000001110010010100;
        11'd1285: TDATA = 37'b0001111011000110011100101110010010001;
        11'd1286: TDATA = 37'b0001111011100011000000101110010001110;
        11'd1287: TDATA = 37'b0001111011111111100011101110010001011;
        11'd1288: TDATA = 37'b0001111100011100000110001110010001000;
        11'd1289: TDATA = 37'b0001111100111000100111101110010000110;
        11'd1290: TDATA = 37'b0001111101010101001000101110010000011;
        11'd1291: TDATA = 37'b0001111101110001101001001110010000000;
        11'd1292: TDATA = 37'b0001111110001110001000101110001111101;
        11'd1293: TDATA = 37'b0001111110101010100111101110001111010;
        11'd1294: TDATA = 37'b0001111111000111000101101110001110111;
        11'd1295: TDATA = 37'b0001111111100011100011001110001110101;
        11'd1296: TDATA = 37'b0010000000000000000000001110001110010;
        11'd1297: TDATA = 37'b0010000000011100011100001110001101111;
        11'd1298: TDATA = 37'b0010000000111000110111101110001101100;
        11'd1299: TDATA = 37'b0010000001010101010010001110001101001;
        11'd1300: TDATA = 37'b0010000001110001101100001110001100111;
        11'd1301: TDATA = 37'b0010000010001110000101101110001100100;
        11'd1302: TDATA = 37'b0010000010101010011110001110001100001;
        11'd1303: TDATA = 37'b0010000011000110110110001110001011110;
        11'd1304: TDATA = 37'b0010000011100011001101001110001011011;
        11'd1305: TDATA = 37'b0010000011111111100011101110001011001;
        11'd1306: TDATA = 37'b0010000100011011111001101110001010110;
        11'd1307: TDATA = 37'b0010000100111000001110101110001010011;
        11'd1308: TDATA = 37'b0010000101010100100011001110001010000;
        11'd1309: TDATA = 37'b0010000101110000110110101110001001110;
        11'd1310: TDATA = 37'b0010000110001101001010001110001001011;
        11'd1311: TDATA = 37'b0010000110101001011100001110001001000;
        11'd1312: TDATA = 37'b0010000111000101101110001110001000101;
        11'd1313: TDATA = 37'b0010000111100001111110101110001000010;
        11'd1314: TDATA = 37'b0010000111111110001111001110001000000;
        11'd1315: TDATA = 37'b0010001000011010011110101110000111101;
        11'd1316: TDATA = 37'b0010001000110110101101101110000111010;
        11'd1317: TDATA = 37'b0010001001010010111011101110000110111;
        11'd1318: TDATA = 37'b0010001001101111001001001110000110101;
        11'd1319: TDATA = 37'b0010001010001011010110001110000110010;
        11'd1320: TDATA = 37'b0010001010100111100010001110000101111;
        11'd1321: TDATA = 37'b0010001011000011101101101110000101101;
        11'd1322: TDATA = 37'b0010001011011111111000101110000101010;
        11'd1323: TDATA = 37'b0010001011111100000010101110000100111;
        11'd1324: TDATA = 37'b0010001100011000001100001110000100100;
        11'd1325: TDATA = 37'b0010001100110100010101001110000100010;
        11'd1326: TDATA = 37'b0010001101010000011101001110000011111;
        11'd1327: TDATA = 37'b0010001101101100100100101110000011100;
        11'd1328: TDATA = 37'b0010001110001000101011001110000011010;
        11'd1329: TDATA = 37'b0010001110100100110001001110000010111;
        11'd1330: TDATA = 37'b0010001111000000110110101110000010100;
        11'd1331: TDATA = 37'b0010001111011100111011001110000010001;
        11'd1332: TDATA = 37'b0010001111111000111111001110000001111;
        11'd1333: TDATA = 37'b0010010000010101000010101110000001100;
        11'd1334: TDATA = 37'b0010010000110001000101001110000001001;
        11'd1335: TDATA = 37'b0010010001001101000111001110000000111;
        11'd1336: TDATA = 37'b0010010001101001001000101110000000100;
        11'd1337: TDATA = 37'b0010010010000101001001001110000000001;
        11'd1338: TDATA = 37'b0010010010100001001001001101111111111;
        11'd1339: TDATA = 37'b0010010010111101001000101101111111100;
        11'd1340: TDATA = 37'b0010010011011001000111001101111111001;
        11'd1341: TDATA = 37'b0010010011110101000101001101111110111;
        11'd1342: TDATA = 37'b0010010100010001000010101101111110100;
        11'd1343: TDATA = 37'b0010010100101100111111001101111110001;
        11'd1344: TDATA = 37'b0010010101001000111011001101111101111;
        11'd1345: TDATA = 37'b0010010101100100110110001101111101100;
        11'd1346: TDATA = 37'b0010010110000000110001001101111101001;
        11'd1347: TDATA = 37'b0010010110011100101011001101111100111;
        11'd1348: TDATA = 37'b0010010110111000100100001101111100100;
        11'd1349: TDATA = 37'b0010010111010100011101001101111100001;
        11'd1350: TDATA = 37'b0010010111110000010101001101111011111;
        11'd1351: TDATA = 37'b0010011000001100001100001101111011100;
        11'd1352: TDATA = 37'b0010011000101000000011001101111011001;
        11'd1353: TDATA = 37'b0010011001000011111001001101111010111;
        11'd1354: TDATA = 37'b0010011001011111101110001101111010100;
        11'd1355: TDATA = 37'b0010011001111011100011001101111010001;
        11'd1356: TDATA = 37'b0010011010010111010111001101111001111;
        11'd1357: TDATA = 37'b0010011010110011001010101101111001100;
        11'd1358: TDATA = 37'b0010011011001110111101001101111001010;
        11'd1359: TDATA = 37'b0010011011101010101111001101111000111;
        11'd1360: TDATA = 37'b0010011100000110100000101101111000100;
        11'd1361: TDATA = 37'b0010011100100010010001101101111000010;
        11'd1362: TDATA = 37'b0010011100111110000001101101110111111;
        11'd1363: TDATA = 37'b0010011101011001110001001101110111101;
        11'd1364: TDATA = 37'b0010011101110101011111101101110111010;
        11'd1365: TDATA = 37'b0010011110010001001110001101110110111;
        11'd1366: TDATA = 37'b0010011110101100111011101101110110101;
        11'd1367: TDATA = 37'b0010011111001000101000001101110110010;
        11'd1368: TDATA = 37'b0010011111100100010100101101110110000;
        11'd1369: TDATA = 37'b0010100000000000000000001101110101101;
        11'd1370: TDATA = 37'b0010100000011011101011001101110101010;
        11'd1371: TDATA = 37'b0010100000110111010101001101110101000;
        11'd1372: TDATA = 37'b0010100001010010111111001101110100101;
        11'd1373: TDATA = 37'b0010100001101110101000001101110100011;
        11'd1374: TDATA = 37'b0010100010001010010000001101110100000;
        11'd1375: TDATA = 37'b0010100010100101111000001101110011101;
        11'd1376: TDATA = 37'b0010100011000001011111001101110011011;
        11'd1377: TDATA = 37'b0010100011011101000101101101110011000;
        11'd1378: TDATA = 37'b0010100011111000101011001101110010110;
        11'd1379: TDATA = 37'b0010100100010100010000001101110010011;
        11'd1380: TDATA = 37'b0010100100101111110100101101110010001;
        11'd1381: TDATA = 37'b0010100101001011011000101101110001110;
        11'd1382: TDATA = 37'b0010100101100110111100001101110001100;
        11'd1383: TDATA = 37'b0010100110000010011110101101110001001;
        11'd1384: TDATA = 37'b0010100110011110000000101101110000110;
        11'd1385: TDATA = 37'b0010100110111001100001101101110000100;
        11'd1386: TDATA = 37'b0010100111010101000010001101110000001;
        11'd1387: TDATA = 37'b0010100111110000100010101101101111111;
        11'd1388: TDATA = 37'b0010101000001100000001101101101111100;
        11'd1389: TDATA = 37'b0010101000100111100000101101101111010;
        11'd1390: TDATA = 37'b0010101001000010111110101101101110111;
        11'd1391: TDATA = 37'b0010101001011110011100001101101110101;
        11'd1392: TDATA = 37'b0010101001111001111001001101101110010;
        11'd1393: TDATA = 37'b0010101010010101010101001101101110000;
        11'd1394: TDATA = 37'b0010101010110000110000101101101101101;
        11'd1395: TDATA = 37'b0010101011001100001011101101101101011;
        11'd1396: TDATA = 37'b0010101011100111100110001101101101000;
        11'd1397: TDATA = 37'b0010101100000011000000001101101100110;
        11'd1398: TDATA = 37'b0010101100011110011001001101101100011;
        11'd1399: TDATA = 37'b0010101100111001110001101101101100001;
        11'd1400: TDATA = 37'b0010101101010101001001001101101011110;
        11'd1401: TDATA = 37'b0010101101110000100000101101101011100;
        11'd1402: TDATA = 37'b0010101110001011110111001101101011001;
        11'd1403: TDATA = 37'b0010101110100111001101001101101010111;
        11'd1404: TDATA = 37'b0010101111000010100010101101101010100;
        11'd1405: TDATA = 37'b0010101111011101110111001101101010010;
        11'd1406: TDATA = 37'b0010101111111001001011001101101001111;
        11'd1407: TDATA = 37'b0010110000010100011110101101101001101;
        11'd1408: TDATA = 37'b0010110000101111110001101101101001010;
        11'd1409: TDATA = 37'b0010110001001011000011101101101001000;
        11'd1410: TDATA = 37'b0010110001100110010101001101101000101;
        11'd1411: TDATA = 37'b0010110010000001100110001101101000011;
        11'd1412: TDATA = 37'b0010110010011100110110101101101000000;
        11'd1413: TDATA = 37'b0010110010111000000110101101100111110;
        11'd1414: TDATA = 37'b0010110011010011010101101101100111011;
        11'd1415: TDATA = 37'b0010110011101110100100001101100111001;
        11'd1416: TDATA = 37'b0010110100001001110010001101100110110;
        11'd1417: TDATA = 37'b0010110100100100111111001101100110100;
        11'd1418: TDATA = 37'b0010110101000000001100001101100110001;
        11'd1419: TDATA = 37'b0010110101011011011000001101100101111;
        11'd1420: TDATA = 37'b0010110101110110100011101101100101101;
        11'd1421: TDATA = 37'b0010110110010001101110101101100101010;
        11'd1422: TDATA = 37'b0010110110101100111000101101100101000;
        11'd1423: TDATA = 37'b0010110111001000000010001101100100101;
        11'd1424: TDATA = 37'b0010110111100011001011001101100100011;
        11'd1425: TDATA = 37'b0010110111111110010011101101100100000;
        11'd1426: TDATA = 37'b0010111000011001011011101101100011110;
        11'd1427: TDATA = 37'b0010111000110100100010101101100011011;
        11'd1428: TDATA = 37'b0010111001001111101001001101100011001;
        11'd1429: TDATA = 37'b0010111001101010101111001101100010111;
        11'd1430: TDATA = 37'b0010111010000101110100101101100010100;
        11'd1431: TDATA = 37'b0010111010100000111001001101100010010;
        11'd1432: TDATA = 37'b0010111010111011111101001101100001111;
        11'd1433: TDATA = 37'b0010111011010111000001001101100001101;
        11'd1434: TDATA = 37'b0010111011110010000011101101100001011;
        11'd1435: TDATA = 37'b0010111100001101000110001101100001000;
        11'd1436: TDATA = 37'b0010111100101000001000001101100000110;
        11'd1437: TDATA = 37'b0010111101000011001001001101100000011;
        11'd1438: TDATA = 37'b0010111101011110001001101101100000001;
        11'd1439: TDATA = 37'b0010111101111001001001101101011111111;
        11'd1440: TDATA = 37'b0010111110010100001000101101011111100;
        11'd1441: TDATA = 37'b0010111110101111000111101101011111010;
        11'd1442: TDATA = 37'b0010111111001010000101101101011110111;
        11'd1443: TDATA = 37'b0010111111100101000011001101011110101;
        11'd1444: TDATA = 37'b0011000000000000000000001101011110011;
        11'd1445: TDATA = 37'b0011000000011010111100101101011110000;
        11'd1446: TDATA = 37'b0011000000110101111000001101011101110;
        11'd1447: TDATA = 37'b0011000001010000110011001101011101011;
        11'd1448: TDATA = 37'b0011000001101011101110001101011101001;
        11'd1449: TDATA = 37'b0011000010000110100111101101011100111;
        11'd1450: TDATA = 37'b0011000010100001100001001101011100100;
        11'd1451: TDATA = 37'b0011000010111100011010001101011100010;
        11'd1452: TDATA = 37'b0011000011010111010010001101011011111;
        11'd1453: TDATA = 37'b0011000011110010001001101101011011101;
        11'd1454: TDATA = 37'b0011000100001101000000101101011011011;
        11'd1455: TDATA = 37'b0011000100100111110111001101011011000;
        11'd1456: TDATA = 37'b0011000101000010101101001101011010110;
        11'd1457: TDATA = 37'b0011000101011101100010001101011010100;
        11'd1458: TDATA = 37'b0011000101111000010110101101011010001;
        11'd1459: TDATA = 37'b0011000110010011001010101101011001111;
        11'd1460: TDATA = 37'b0011000110101101111110001101011001101;
        11'd1461: TDATA = 37'b0011000111001000110001001101011001010;
        11'd1462: TDATA = 37'b0011000111100011100011001101011001000;
        11'd1463: TDATA = 37'b0011000111111110010101001101011000110;
        11'd1464: TDATA = 37'b0011001000011001000110001101011000011;
        11'd1465: TDATA = 37'b0011001000110011110110101101011000001;
        11'd1466: TDATA = 37'b0011001001001110100110101101010111111;
        11'd1467: TDATA = 37'b0011001001101001010110001101010111100;
        11'd1468: TDATA = 37'b0011001010000100000100101101010111010;
        11'd1469: TDATA = 37'b0011001010011110110011001101010111000;
        11'd1470: TDATA = 37'b0011001010111001100000101101010110101;
        11'd1471: TDATA = 37'b0011001011010100001101101101010110011;
        11'd1472: TDATA = 37'b0011001011101110111010001101010110001;
        11'd1473: TDATA = 37'b0011001100001001100101101101010101110;
        11'd1474: TDATA = 37'b0011001100100100010001001101010101100;
        11'd1475: TDATA = 37'b0011001100111110111011101101010101010;
        11'd1476: TDATA = 37'b0011001101011001100110001101010100111;
        11'd1477: TDATA = 37'b0011001101110100001111101101010100101;
        11'd1478: TDATA = 37'b0011001110001110111000101101010100011;
        11'd1479: TDATA = 37'b0011001110101001100000101101010100000;
        11'd1480: TDATA = 37'b0011001111000100001000101101010011110;
        11'd1481: TDATA = 37'b0011001111011110110000001101010011100;
        11'd1482: TDATA = 37'b0011001111111001010110101101010011010;
        11'd1483: TDATA = 37'b0011010000010011111100101101010010111;
        11'd1484: TDATA = 37'b0011010000101110100010001101010010101;
        11'd1485: TDATA = 37'b0011010001001001000111001101010010011;
        11'd1486: TDATA = 37'b0011010001100011101011101101010010000;
        11'd1487: TDATA = 37'b0011010001111110001111001101010001110;
        11'd1488: TDATA = 37'b0011010010011000110010101101010001100;
        11'd1489: TDATA = 37'b0011010010110011010101001101010001001;
        11'd1490: TDATA = 37'b0011010011001101110111001101010000111;
        11'd1491: TDATA = 37'b0011010011101000011000101101010000101;
        11'd1492: TDATA = 37'b0011010100000010111001101101010000011;
        11'd1493: TDATA = 37'b0011010100011101011010001101010000000;
        11'd1494: TDATA = 37'b0011010100110111111010001101001111110;
        11'd1495: TDATA = 37'b0011010101010010011001001101001111100;
        11'd1496: TDATA = 37'b0011010101101100110111101101001111010;
        11'd1497: TDATA = 37'b0011010110000111010110001101001110111;
        11'd1498: TDATA = 37'b0011010110100001110011101101001110101;
        11'd1499: TDATA = 37'b0011010110111100010000101101001110011;
        11'd1500: TDATA = 37'b0011010111010110101100101101001110001;
        11'd1501: TDATA = 37'b0011010111110001001000101101001101110;
        11'd1502: TDATA = 37'b0011011000001011100100001101001101100;
        11'd1503: TDATA = 37'b0011011000100101111110101101001101010;
        11'd1504: TDATA = 37'b0011011001000000011001001101001101000;
        11'd1505: TDATA = 37'b0011011001011010110010101101001100101;
        11'd1506: TDATA = 37'b0011011001110101001011101101001100011;
        11'd1507: TDATA = 37'b0011011010001111100100001101001100001;
        11'd1508: TDATA = 37'b0011011010101001111100001101001011111;
        11'd1509: TDATA = 37'b0011011011000100010011001101001011100;
        11'd1510: TDATA = 37'b0011011011011110101010001101001011010;
        11'd1511: TDATA = 37'b0011011011111001000000001101001011000;
        11'd1512: TDATA = 37'b0011011100010011010110001101001010110;
        11'd1513: TDATA = 37'b0011011100101101101011001101001010011;
        11'd1514: TDATA = 37'b0011011101000111111111101101001010001;
        11'd1515: TDATA = 37'b0011011101100010010011101101001001111;
        11'd1516: TDATA = 37'b0011011101111100100111001101001001101;
        11'd1517: TDATA = 37'b0011011110010110111010001101001001010;
        11'd1518: TDATA = 37'b0011011110110001001100101101001001000;
        11'd1519: TDATA = 37'b0011011111001011011110001101001000110;
        11'd1520: TDATA = 37'b0011011111100101101111101101001000100;
        11'd1521: TDATA = 37'b0011100000000000000000001101001000010;
        11'd1522: TDATA = 37'b0011100000011010010000001101000111111;
        11'd1523: TDATA = 37'b0011100000110100011111101101000111101;
        11'd1524: TDATA = 37'b0011100001001110101110101101000111011;
        11'd1525: TDATA = 37'b0011100001101000111101001101000111001;
        11'd1526: TDATA = 37'b0011100010000011001011001101000110111;
        11'd1527: TDATA = 37'b0011100010011101011000101101000110100;
        11'd1528: TDATA = 37'b0011100010110111100101101101000110010;
        11'd1529: TDATA = 37'b0011100011010001110001101101000110000;
        11'd1530: TDATA = 37'b0011100011101011111101101101000101110;
        11'd1531: TDATA = 37'b0011100100000110001000101101000101100;
        11'd1532: TDATA = 37'b0011100100100000010011001101000101001;
        11'd1533: TDATA = 37'b0011100100111010011101101101000100111;
        11'd1534: TDATA = 37'b0011100101010100100111001101000100101;
        11'd1535: TDATA = 37'b0011100101101110110000001101000100011;
        11'd1536: TDATA = 37'b0011100110001000111000101101000100001;
        11'd1537: TDATA = 37'b0011100110100011000000001101000011111;
        11'd1538: TDATA = 37'b0011100110111101000111101101000011100;
        11'd1539: TDATA = 37'b0011100111010111001110101101000011010;
        11'd1540: TDATA = 37'b0011100111110001010100101101000011000;
        11'd1541: TDATA = 37'b0011101000001011011010101101000010110;
        11'd1542: TDATA = 37'b0011101000100101011111101101000010100;
        11'd1543: TDATA = 37'b0011101000111111100100101101000010010;
        11'd1544: TDATA = 37'b0011101001011001101000101101000001111;
        11'd1545: TDATA = 37'b0011101001110011101100001101000001101;
        11'd1546: TDATA = 37'b0011101010001101101111001101000001011;
        11'd1547: TDATA = 37'b0011101010100111110001101101000001001;
        11'd1548: TDATA = 37'b0011101011000001110011101101000000111;
        11'd1549: TDATA = 37'b0011101011011011110101001101000000101;
        11'd1550: TDATA = 37'b0011101011110101110110001101000000010;
        11'd1551: TDATA = 37'b0011101100001111110110001101000000000;
        11'd1552: TDATA = 37'b0011101100101001110110001100111111110;
        11'd1553: TDATA = 37'b0011101101000011110101001100111111100;
        11'd1554: TDATA = 37'b0011101101011101110100001100111111010;
        11'd1555: TDATA = 37'b0011101101110111110010001100111111000;
        11'd1556: TDATA = 37'b0011101110010001110000001100111110110;
        11'd1557: TDATA = 37'b0011101110101011101101001100111110011;
        11'd1558: TDATA = 37'b0011101111000101101001101100111110001;
        11'd1559: TDATA = 37'b0011101111011111100101101100111101111;
        11'd1560: TDATA = 37'b0011101111111001100001001100111101101;
        11'd1561: TDATA = 37'b0011110000010011011100001100111101011;
        11'd1562: TDATA = 37'b0011110000101101010110101100111101001;
        11'd1563: TDATA = 37'b0011110001000111010000101100111100111;
        11'd1564: TDATA = 37'b0011110001100001001010001100111100101;
        11'd1565: TDATA = 37'b0011110001111011000011001100111100010;
        11'd1566: TDATA = 37'b0011110010010100111011101100111100000;
        11'd1567: TDATA = 37'b0011110010101110110011001100111011110;
        11'd1568: TDATA = 37'b0011110011001000101010101100111011100;
        11'd1569: TDATA = 37'b0011110011100010100001001100111011010;
        11'd1570: TDATA = 37'b0011110011111100010111101100111011000;
        11'd1571: TDATA = 37'b0011110100010110001101001100111010110;
        11'd1572: TDATA = 37'b0011110100110000000010101100111010100;
        11'd1573: TDATA = 37'b0011110101001001110111001100111010010;
        11'd1574: TDATA = 37'b0011110101100011101011001100111010000;
        11'd1575: TDATA = 37'b0011110101111101011110101100111001101;
        11'd1576: TDATA = 37'b0011110110010111010010001100111001011;
        11'd1577: TDATA = 37'b0011110110110001000100101100111001001;
        11'd1578: TDATA = 37'b0011110111001010110110101100111000111;
        11'd1579: TDATA = 37'b0011110111100100101000001100111000101;
        11'd1580: TDATA = 37'b0011110111111110011001001100111000011;
        11'd1581: TDATA = 37'b0011111000011000001001101100111000001;
        11'd1582: TDATA = 37'b0011111000110001111001101100110111111;
        11'd1583: TDATA = 37'b0011111001001011101001001100110111101;
        11'd1584: TDATA = 37'b0011111001100101010111101100110111011;
        11'd1585: TDATA = 37'b0011111001111111000110001100110111001;
        11'd1586: TDATA = 37'b0011111010011000110100001100110110110;
        11'd1587: TDATA = 37'b0011111010110010100001101100110110100;
        11'd1588: TDATA = 37'b0011111011001100001110001100110110010;
        11'd1589: TDATA = 37'b0011111011100101111010101100110110000;
        11'd1590: TDATA = 37'b0011111011111111100110101100110101110;
        11'd1591: TDATA = 37'b0011111100011001010001101100110101100;
        11'd1592: TDATA = 37'b0011111100110010111100101100110101010;
        11'd1593: TDATA = 37'b0011111101001100100110101100110101000;
        11'd1594: TDATA = 37'b0011111101100110010000101100110100110;
        11'd1595: TDATA = 37'b0011111101111111111001101100110100100;
        11'd1596: TDATA = 37'b0011111110011001100010101100110100010;
        11'd1597: TDATA = 37'b0011111110110011001010101100110100000;
        11'd1598: TDATA = 37'b0011111111001100110010001100110011110;
        11'd1599: TDATA = 37'b0011111111100110011001101100110011100;
        11'd1600: TDATA = 37'b0100000000000000000000001100110011010;
        11'd1601: TDATA = 37'b0100000000011001100110001100110011000;
        11'd1602: TDATA = 37'b0100000000110011001100001100110010110;
        11'd1603: TDATA = 37'b0100000001001100110001001100110010011;
        11'd1604: TDATA = 37'b0100000001100110010101101100110010001;
        11'd1605: TDATA = 37'b0100000001111111111001101100110001111;
        11'd1606: TDATA = 37'b0100000010011001011101001100110001101;
        11'd1607: TDATA = 37'b0100000010110011000000101100110001011;
        11'd1608: TDATA = 37'b0100000011001100100011001100110001001;
        11'd1609: TDATA = 37'b0100000011100110000101001100110000111;
        11'd1610: TDATA = 37'b0100000011111111100110101100110000101;
        11'd1611: TDATA = 37'b0100000100011001000111101100110000011;
        11'd1612: TDATA = 37'b0100000100110010101000001100110000001;
        11'd1613: TDATA = 37'b0100000101001100001000001100101111111;
        11'd1614: TDATA = 37'b0100000101100101100111101100101111101;
        11'd1615: TDATA = 37'b0100000101111111000110101100101111011;
        11'd1616: TDATA = 37'b0100000110011000100101001100101111001;
        11'd1617: TDATA = 37'b0100000110110010000011001100101110111;
        11'd1618: TDATA = 37'b0100000111001011100000101100101110101;
        11'd1619: TDATA = 37'b0100000111100100111101101100101110011;
        11'd1620: TDATA = 37'b0100000111111110011010001100101110001;
        11'd1621: TDATA = 37'b0100001000010111110110001100101101111;
        11'd1622: TDATA = 37'b0100001000110001010001101100101101101;
        11'd1623: TDATA = 37'b0100001001001010101100101100101101011;
        11'd1624: TDATA = 37'b0100001001100100000111001100101101001;
        11'd1625: TDATA = 37'b0100001001111101100001001100101100111;
        11'd1626: TDATA = 37'b0100001010010110111010101100101100101;
        11'd1627: TDATA = 37'b0100001010110000010011101100101100011;
        11'd1628: TDATA = 37'b0100001011001001101100001100101100001;
        11'd1629: TDATA = 37'b0100001011100011000100001100101011111;
        11'd1630: TDATA = 37'b0100001011111100011011101100101011101;
        11'd1631: TDATA = 37'b0100001100010101110010101100101011011;
        11'd1632: TDATA = 37'b0100001100101111001001001100101011001;
        11'd1633: TDATA = 37'b0100001101001000011111101100101010111;
        11'd1634: TDATA = 37'b0100001101100001110101001100101010101;
        11'd1635: TDATA = 37'b0100001101111011001010001100101010011;
        11'd1636: TDATA = 37'b0100001110010100011110101100101010001;
        11'd1637: TDATA = 37'b0100001110101101110010101100101001111;
        11'd1638: TDATA = 37'b0100001111000111000110001100101001101;
        11'd1639: TDATA = 37'b0100001111100000011001001100101001011;
        11'd1640: TDATA = 37'b0100001111111001101011101100101001001;
        11'd1641: TDATA = 37'b0100010000010010111101101100101000111;
        11'd1642: TDATA = 37'b0100010000101100001111001100101000101;
        11'd1643: TDATA = 37'b0100010001000101100000001100101000011;
        11'd1644: TDATA = 37'b0100010001011110110000101100101000001;
        11'd1645: TDATA = 37'b0100010001111000000001001100100111111;
        11'd1646: TDATA = 37'b0100010010010001010000101100100111101;
        11'd1647: TDATA = 37'b0100010010101010011111101100100111011;
        11'd1648: TDATA = 37'b0100010011000011101110001100100111001;
        11'd1649: TDATA = 37'b0100010011011100111100001100100110111;
        11'd1650: TDATA = 37'b0100010011110110001010001100100110110;
        11'd1651: TDATA = 37'b0100010100001111010111001100100110100;
        11'd1652: TDATA = 37'b0100010100101000100011101100100110010;
        11'd1653: TDATA = 37'b0100010101000001110000001100100110000;
        11'd1654: TDATA = 37'b0100010101011010111011101100100101110;
        11'd1655: TDATA = 37'b0100010101110100000110101100100101100;
        11'd1656: TDATA = 37'b0100010110001101010001101100100101010;
        11'd1657: TDATA = 37'b0100010110100110011011101100100101000;
        11'd1658: TDATA = 37'b0100010110111111100101101100100100110;
        11'd1659: TDATA = 37'b0100010111011000101110101100100100100;
        11'd1660: TDATA = 37'b0100010111110001110111101100100100010;
        11'd1661: TDATA = 37'b0100011000001010111111101100100100000;
        11'd1662: TDATA = 37'b0100011000100100000111101100100011110;
        11'd1663: TDATA = 37'b0100011000111101001110101100100011100;
        11'd1664: TDATA = 37'b0100011001010110010101101100100011010;
        11'd1665: TDATA = 37'b0100011001101111011100001100100011000;
        11'd1666: TDATA = 37'b0100011010001000100001101100100010110;
        11'd1667: TDATA = 37'b0100011010100001100111001100100010101;
        11'd1668: TDATA = 37'b0100011010111010101100001100100010011;
        11'd1669: TDATA = 37'b0100011011010011110000101100100010001;
        11'd1670: TDATA = 37'b0100011011101100110100101100100001111;
        11'd1671: TDATA = 37'b0100011100000101111000001100100001101;
        11'd1672: TDATA = 37'b0100011100011110111010101100100001011;
        11'd1673: TDATA = 37'b0100011100110111111101001100100001001;
        11'd1674: TDATA = 37'b0100011101010000111111101100100000111;
        11'd1675: TDATA = 37'b0100011101101010000001001100100000101;
        11'd1676: TDATA = 37'b0100011110000011000010001100100000011;
        11'd1677: TDATA = 37'b0100011110011100000010101100100000001;
        11'd1678: TDATA = 37'b0100011110110101000010101100011111111;
        11'd1679: TDATA = 37'b0100011111001110000010001100011111110;
        11'd1680: TDATA = 37'b0100011111100111000001101100011111100;
        11'd1681: TDATA = 37'b0100100000000000000000001100011111010;
        11'd1682: TDATA = 37'b0100100000011000111110001100011111000;
        11'd1683: TDATA = 37'b0100100000110001111100001100011110110;
        11'd1684: TDATA = 37'b0100100001001010111001001100011110100;
        11'd1685: TDATA = 37'b0100100001100011110110001100011110010;
        11'd1686: TDATA = 37'b0100100001111100110010101100011110000;
        11'd1687: TDATA = 37'b0100100010010101101110001100011101110;
        11'd1688: TDATA = 37'b0100100010101110101001101100011101100;
        11'd1689: TDATA = 37'b0100100011000111100100101100011101011;
        11'd1690: TDATA = 37'b0100100011100000011110101100011101001;
        11'd1691: TDATA = 37'b0100100011111001011000101100011100111;
        11'd1692: TDATA = 37'b0100100100010010010010001100011100101;
        11'd1693: TDATA = 37'b0100100100101011001011001100011100011;
        11'd1694: TDATA = 37'b0100100101000100000011101100011100001;
        11'd1695: TDATA = 37'b0100100101011100111011101100011011111;
        11'd1696: TDATA = 37'b0100100101110101110011101100011011101;
        11'd1697: TDATA = 37'b0100100110001110101010101100011011100;
        11'd1698: TDATA = 37'b0100100110100111100001001100011011010;
        11'd1699: TDATA = 37'b0100100111000000010111101100011011000;
        11'd1700: TDATA = 37'b0100100111011001001101001100011010110;
        11'd1701: TDATA = 37'b0100100111110010000010101100011010100;
        11'd1702: TDATA = 37'b0100101000001010110111001100011010010;
        11'd1703: TDATA = 37'b0100101000100011101011101100011010000;
        11'd1704: TDATA = 37'b0100101000111100011111001100011001110;
        11'd1705: TDATA = 37'b0100101001010101010010101100011001101;
        11'd1706: TDATA = 37'b0100101001101110000101101100011001011;
        11'd1707: TDATA = 37'b0100101010000110111000001100011001001;
        11'd1708: TDATA = 37'b0100101010011111101010001100011000111;
        11'd1709: TDATA = 37'b0100101010111000011011101100011000101;
        11'd1710: TDATA = 37'b0100101011010001001100101100011000011;
        11'd1711: TDATA = 37'b0100101011101001111101001100011000001;
        11'd1712: TDATA = 37'b0100101100000010101101001100011000000;
        11'd1713: TDATA = 37'b0100101100011011011101001100010111110;
        11'd1714: TDATA = 37'b0100101100110100001100001100010111100;
        11'd1715: TDATA = 37'b0100101101001100111011001100010111010;
        11'd1716: TDATA = 37'b0100101101100101101001001100010111000;
        11'd1717: TDATA = 37'b0100101101111110010111001100010110110;
        11'd1718: TDATA = 37'b0100101110010111000100101100010110101;
        11'd1719: TDATA = 37'b0100101110101111110001001100010110011;
        11'd1720: TDATA = 37'b0100101111001000011101101100010110001;
        11'd1721: TDATA = 37'b0100101111100001001001101100010101111;
        11'd1722: TDATA = 37'b0100101111111001110101001100010101101;
        11'd1723: TDATA = 37'b0100110000010010100000101100010101011;
        11'd1724: TDATA = 37'b0100110000101011001011001100010101010;
        11'd1725: TDATA = 37'b0100110001000011110101001100010101000;
        11'd1726: TDATA = 37'b0100110001011100011110101100010100110;
        11'd1727: TDATA = 37'b0100110001110101001000001100010100100;
        11'd1728: TDATA = 37'b0100110010001101110000101100010100010;
        11'd1729: TDATA = 37'b0100110010100110011001001100010100000;
        11'd1730: TDATA = 37'b0100110010111111000001001100010011111;
        11'd1731: TDATA = 37'b0100110011010111101000101100010011101;
        11'd1732: TDATA = 37'b0100110011110000001111101100010011011;
        11'd1733: TDATA = 37'b0100110100001000110110001100010011001;
        11'd1734: TDATA = 37'b0100110100100001011100001100010010111;
        11'd1735: TDATA = 37'b0100110100111010000001101100010010101;
        11'd1736: TDATA = 37'b0100110101010010100110101100010010100;
        11'd1737: TDATA = 37'b0100110101101011001011101100010010010;
        11'd1738: TDATA = 37'b0100110110000011101111101100010010000;
        11'd1739: TDATA = 37'b0100110110011100010011101100010001110;
        11'd1740: TDATA = 37'b0100110110110100110110101100010001100;
        11'd1741: TDATA = 37'b0100110111001101011001101100010001011;
        11'd1742: TDATA = 37'b0100110111100101111100001100010001001;
        11'd1743: TDATA = 37'b0100110111111110011110001100010000111;
        11'd1744: TDATA = 37'b0100111000010110111111101100010000101;
        11'd1745: TDATA = 37'b0100111000101111100000101100010000011;
        11'd1746: TDATA = 37'b0100111001001000000001001100010000010;
        11'd1747: TDATA = 37'b0100111001100000100001101100010000000;
        11'd1748: TDATA = 37'b0100111001111001000001001100001111110;
        11'd1749: TDATA = 37'b0100111010010001100000101100001111100;
        11'd1750: TDATA = 37'b0100111010101001111111001100001111010;
        11'd1751: TDATA = 37'b0100111011000010011101101100001111001;
        11'd1752: TDATA = 37'b0100111011011010111011101100001110111;
        11'd1753: TDATA = 37'b0100111011110011011001001100001110101;
        11'd1754: TDATA = 37'b0100111100001011110110001100001110011;
        11'd1755: TDATA = 37'b0100111100100100010010101100001110010;
        11'd1756: TDATA = 37'b0100111100111100101111001100001110000;
        11'd1757: TDATA = 37'b0100111101010101001010101100001101110;
        11'd1758: TDATA = 37'b0100111101101101100101101100001101100;
        11'd1759: TDATA = 37'b0100111110000110000000101100001101010;
        11'd1760: TDATA = 37'b0100111110011110011011001100001101001;
        11'd1761: TDATA = 37'b0100111110110110110101001100001100111;
        11'd1762: TDATA = 37'b0100111111001111001110101100001100101;
        11'd1763: TDATA = 37'b0100111111100111100111101100001100011;
        11'd1764: TDATA = 37'b0101000000000000000000001100001100010;
        11'd1765: TDATA = 37'b0101000000011000011000001100001100000;
        11'd1766: TDATA = 37'b0101000000110000110000001100001011110;
        11'd1767: TDATA = 37'b0101000001001001000111001100001011100;
        11'd1768: TDATA = 37'b0101000001100001011110001100001011010;
        11'd1769: TDATA = 37'b0101000001111001110100101100001011001;
        11'd1770: TDATA = 37'b0101000010010010001010101100001010111;
        11'd1771: TDATA = 37'b0101000010101010100000001100001010101;
        11'd1772: TDATA = 37'b0101000011000010110101001100001010011;
        11'd1773: TDATA = 37'b0101000011011011001001101100001010010;
        11'd1774: TDATA = 37'b0101000011110011011110001100001010000;
        11'd1775: TDATA = 37'b0101000100001011110001101100001001110;
        11'd1776: TDATA = 37'b0101000100100100000101001100001001100;
        11'd1777: TDATA = 37'b0101000100111100010111101100001001011;
        11'd1778: TDATA = 37'b0101000101010100101010001100001001001;
        11'd1779: TDATA = 37'b0101000101101100111100001100001000111;
        11'd1780: TDATA = 37'b0101000110000101001101101100001000101;
        11'd1781: TDATA = 37'b0101000110011101011111001100001000100;
        11'd1782: TDATA = 37'b0101000110110101101111101100001000010;
        11'd1783: TDATA = 37'b0101000111001110000000001100001000000;
        11'd1784: TDATA = 37'b0101000111100110001111101100000111110;
        11'd1785: TDATA = 37'b0101000111111110011111001100000111101;
        11'd1786: TDATA = 37'b0101001000010110101110001100000111011;
        11'd1787: TDATA = 37'b0101001000101110111100101100000111001;
        11'd1788: TDATA = 37'b0101001001000111001010101100000110111;
        11'd1789: TDATA = 37'b0101001001011111011000101100000110110;
        11'd1790: TDATA = 37'b0101001001110111100101101100000110100;
        11'd1791: TDATA = 37'b0101001010001111110010101100000110010;
        11'd1792: TDATA = 37'b0101001010100111111110101100000110001;
        11'd1793: TDATA = 37'b0101001011000000001010101100000101111;
        11'd1794: TDATA = 37'b0101001011011000010110001100000101101;
        11'd1795: TDATA = 37'b0101001011110000100001001100000101011;
        11'd1796: TDATA = 37'b0101001100001000101100001100000101010;
        11'd1797: TDATA = 37'b0101001100100000110110001100000101000;
        11'd1798: TDATA = 37'b0101001100111000111111101100000100110;
        11'd1799: TDATA = 37'b0101001101010001001001001100000100101;
        11'd1800: TDATA = 37'b0101001101101001010010001100000100011;
        11'd1801: TDATA = 37'b0101001110000001011010101100000100001;
        11'd1802: TDATA = 37'b0101001110011001100010101100000011111;
        11'd1803: TDATA = 37'b0101001110110001101010001100000011110;
        11'd1804: TDATA = 37'b0101001111001001110001101100000011100;
        11'd1805: TDATA = 37'b0101001111100001111000001100000011010;
        11'd1806: TDATA = 37'b0101001111111001111110101100000011001;
        11'd1807: TDATA = 37'b0101010000010010000100101100000010111;
        11'd1808: TDATA = 37'b0101010000101010001010001100000010101;
        11'd1809: TDATA = 37'b0101010001000010001111001100000010011;
        11'd1810: TDATA = 37'b0101010001011010010011101100000010010;
        11'd1811: TDATA = 37'b0101010001110010011000001100000010000;
        11'd1812: TDATA = 37'b0101010010001010011011101100000001110;
        11'd1813: TDATA = 37'b0101010010100010011111001100000001101;
        11'd1814: TDATA = 37'b0101010010111010100010001100000001011;
        11'd1815: TDATA = 37'b0101010011010010100100101100000001001;
        11'd1816: TDATA = 37'b0101010011101010100110101100000001000;
        11'd1817: TDATA = 37'b0101010100000010101000001100000000110;
        11'd1818: TDATA = 37'b0101010100011010101001101100000000100;
        11'd1819: TDATA = 37'b0101010100110010101010001100000000010;
        11'd1820: TDATA = 37'b0101010101001010101010101100000000001;
        11'd1821: TDATA = 37'b0101010101100010101010101011111111111;
        11'd1822: TDATA = 37'b0101010101111010101010001011111111101;
        11'd1823: TDATA = 37'b0101010110010010101001101011111111100;
        11'd1824: TDATA = 37'b0101010110101010101000001011111111010;
        11'd1825: TDATA = 37'b0101010111000010100110101011111111000;
        11'd1826: TDATA = 37'b0101010111011010100100001011111110111;
        11'd1827: TDATA = 37'b0101010111110010100001101011111110101;
        11'd1828: TDATA = 37'b0101011000001010011110101011111110011;
        11'd1829: TDATA = 37'b0101011000100010011011101011111110010;
        11'd1830: TDATA = 37'b0101011000111010010111101011111110000;
        11'd1831: TDATA = 37'b0101011001010010010011001011111101110;
        11'd1832: TDATA = 37'b0101011001101010001110101011111101101;
        11'd1833: TDATA = 37'b0101011010000010001001101011111101011;
        11'd1834: TDATA = 37'b0101011010011010000100001011111101001;
        11'd1835: TDATA = 37'b0101011010110001111110001011111101000;
        11'd1836: TDATA = 37'b0101011011001001111000001011111100110;
        11'd1837: TDATA = 37'b0101011011100001110001001011111100100;
        11'd1838: TDATA = 37'b0101011011111001101010001011111100011;
        11'd1839: TDATA = 37'b0101011100010001100010101011111100001;
        11'd1840: TDATA = 37'b0101011100101001011010101011111011111;
        11'd1841: TDATA = 37'b0101011101000001010010001011111011110;
        11'd1842: TDATA = 37'b0101011101011001001001001011111011100;
        11'd1843: TDATA = 37'b0101011101110001000000001011111011010;
        11'd1844: TDATA = 37'b0101011110001000110110101011111011001;
        11'd1845: TDATA = 37'b0101011110100000101100101011111010111;
        11'd1846: TDATA = 37'b0101011110111000100010001011111010101;
        11'd1847: TDATA = 37'b0101011111010000010111001011111010100;
        11'd1848: TDATA = 37'b0101011111101000001011101011111010010;
        11'd1849: TDATA = 37'b0101100000000000000000001011111010000;
        11'd1850: TDATA = 37'b0101100000010111110100001011111001111;
        11'd1851: TDATA = 37'b0101100000101111100111101011111001101;
        11'd1852: TDATA = 37'b0101100001000111011010101011111001011;
        11'd1853: TDATA = 37'b0101100001011111001101001011111001010;
        11'd1854: TDATA = 37'b0101100001110110111111101011111001000;
        11'd1855: TDATA = 37'b0101100010001110110001001011111000111;
        11'd1856: TDATA = 37'b0101100010100110100010101011111000101;
        11'd1857: TDATA = 37'b0101100010111110010011101011111000011;
        11'd1858: TDATA = 37'b0101100011010110000100001011111000010;
        11'd1859: TDATA = 37'b0101100011101101110100101011111000000;
        11'd1860: TDATA = 37'b0101100100000101100100001011110111110;
        11'd1861: TDATA = 37'b0101100100011101010011101011110111101;
        11'd1862: TDATA = 37'b0101100100110101000010101011110111011;
        11'd1863: TDATA = 37'b0101100101001100110001001011110111001;
        11'd1864: TDATA = 37'b0101100101100100011111001011110111000;
        11'd1865: TDATA = 37'b0101100101111100001101001011110110110;
        11'd1866: TDATA = 37'b0101100110010011111010101011110110101;
        11'd1867: TDATA = 37'b0101100110101011100111001011110110011;
        11'd1868: TDATA = 37'b0101100111000011010100001011110110001;
        11'd1869: TDATA = 37'b0101100111011011000000001011110110000;
        11'd1870: TDATA = 37'b0101100111110010101011101011110101110;
        11'd1871: TDATA = 37'b0101101000001010010111001011110101100;
        11'd1872: TDATA = 37'b0101101000100010000010001011110101011;
        11'd1873: TDATA = 37'b0101101000111001101100101011110101001;
        11'd1874: TDATA = 37'b0101101001010001010110101011110101000;
        11'd1875: TDATA = 37'b0101101001101001000000001011110100110;
        11'd1876: TDATA = 37'b0101101010000000101001101011110100100;
        11'd1877: TDATA = 37'b0101101010011000010010101011110100011;
        11'd1878: TDATA = 37'b0101101010101111111010101011110100001;
        11'd1879: TDATA = 37'b0101101011000111100011001011110100000;
        11'd1880: TDATA = 37'b0101101011011111001010101011110011110;
        11'd1881: TDATA = 37'b0101101011110110110010001011110011100;
        11'd1882: TDATA = 37'b0101101100001110011000101011110011011;
        11'd1883: TDATA = 37'b0101101100100101111111001011110011001;
        11'd1884: TDATA = 37'b0101101100111101100101001011110010111;
        11'd1885: TDATA = 37'b0101101101010101001011001011110010110;
        11'd1886: TDATA = 37'b0101101101101100110000001011110010100;
        11'd1887: TDATA = 37'b0101101110000100010101001011110010011;
        11'd1888: TDATA = 37'b0101101110011011111001101011110010001;
        11'd1889: TDATA = 37'b0101101110110011011101101011110001111;
        11'd1890: TDATA = 37'b0101101111001011000001001011110001110;
        11'd1891: TDATA = 37'b0101101111100010100100101011110001100;
        11'd1892: TDATA = 37'b0101101111111010000111101011110001011;
        11'd1893: TDATA = 37'b0101110000010001101010001011110001001;
        11'd1894: TDATA = 37'b0101110000101001001100001011110001000;
        11'd1895: TDATA = 37'b0101110001000000101101101011110000110;
        11'd1896: TDATA = 37'b0101110001011000001111001011110000100;
        11'd1897: TDATA = 37'b0101110001101111101111101011110000011;
        11'd1898: TDATA = 37'b0101110010000111010000001011110000001;
        11'd1899: TDATA = 37'b0101110010011110110000101011110000000;
        11'd1900: TDATA = 37'b0101110010110110010000001011101111110;
        11'd1901: TDATA = 37'b0101110011001101101111101011101111100;
        11'd1902: TDATA = 37'b0101110011100101001110001011101111011;
        11'd1903: TDATA = 37'b0101110011111100101100101011101111001;
        11'd1904: TDATA = 37'b0101110100010100001011001011101111000;
        11'd1905: TDATA = 37'b0101110100101011101000101011101110110;
        11'd1906: TDATA = 37'b0101110101000011000110001011101110101;
        11'd1907: TDATA = 37'b0101110101011010100011001011101110011;
        11'd1908: TDATA = 37'b0101110101110001111111101011101110001;
        11'd1909: TDATA = 37'b0101110110001001011011101011101110000;
        11'd1910: TDATA = 37'b0101110110100000110111101011101101110;
        11'd1911: TDATA = 37'b0101110110111000010010101011101101101;
        11'd1912: TDATA = 37'b0101110111001111101101101011101101011;
        11'd1913: TDATA = 37'b0101110111100111001000001011101101010;
        11'd1914: TDATA = 37'b0101110111111110100010101011101101000;
        11'd1915: TDATA = 37'b0101111000010101111100001011101100110;
        11'd1916: TDATA = 37'b0101111000101101010101101011101100101;
        11'd1917: TDATA = 37'b0101111001000100101110101011101100011;
        11'd1918: TDATA = 37'b0101111001011100000111001011101100010;
        11'd1919: TDATA = 37'b0101111001110011011111101011101100000;
        11'd1920: TDATA = 37'b0101111010001010110111101011101011111;
        11'd1921: TDATA = 37'b0101111010100010001110101011101011101;
        11'd1922: TDATA = 37'b0101111010111001100110001011101011011;
        11'd1923: TDATA = 37'b0101111011010000111100101011101011010;
        11'd1924: TDATA = 37'b0101111011101000010011001011101011000;
        11'd1925: TDATA = 37'b0101111011111111101000101011101010111;
        11'd1926: TDATA = 37'b0101111100010110111110001011101010101;
        11'd1927: TDATA = 37'b0101111100101110010011101011101010100;
        11'd1928: TDATA = 37'b0101111101000101101000001011101010010;
        11'd1929: TDATA = 37'b0101111101011100111100101011101010001;
        11'd1930: TDATA = 37'b0101111101110100010000101011101001111;
        11'd1931: TDATA = 37'b0101111110001011100100001011101001110;
        11'd1932: TDATA = 37'b0101111110100010110111001011101001100;
        11'd1933: TDATA = 37'b0101111110111010001010001011101001010;
        11'd1934: TDATA = 37'b0101111111010001011100101011101001001;
        11'd1935: TDATA = 37'b0101111111101000101110101011101000111;
        11'd1936: TDATA = 37'b0110000000000000000000001011101000110;
        11'd1937: TDATA = 37'b0110000000010111010001101011101000100;
        11'd1938: TDATA = 37'b0110000000101110100010001011101000011;
        11'd1939: TDATA = 37'b0110000001000101110010101011101000001;
        11'd1940: TDATA = 37'b0110000001011101000010101011101000000;
        11'd1941: TDATA = 37'b0110000001110100010010101011100111110;
        11'd1942: TDATA = 37'b0110000010001011100010001011100111101;
        11'd1943: TDATA = 37'b0110000010100010110001001011100111011;
        11'd1944: TDATA = 37'b0110000010111001111111101011100111010;
        11'd1945: TDATA = 37'b0110000011010001001101101011100111000;
        11'd1946: TDATA = 37'b0110000011101000011011101011100110110;
        11'd1947: TDATA = 37'b0110000011111111101001001011100110101;
        11'd1948: TDATA = 37'b0110000100010110110110001011100110011;
        11'd1949: TDATA = 37'b0110000100101110000010101011100110010;
        11'd1950: TDATA = 37'b0110000101000101001111001011100110000;
        11'd1951: TDATA = 37'b0110000101011100011010101011100101111;
        11'd1952: TDATA = 37'b0110000101110011100110001011100101101;
        11'd1953: TDATA = 37'b0110000110001010110001101011100101100;
        11'd1954: TDATA = 37'b0110000110100001111100001011100101010;
        11'd1955: TDATA = 37'b0110000110111001000110101011100101001;
        11'd1956: TDATA = 37'b0110000111010000010000101011100100111;
        11'd1957: TDATA = 37'b0110000111100111011010001011100100110;
        11'd1958: TDATA = 37'b0110000111111110100011101011100100100;
        11'd1959: TDATA = 37'b0110001000010101101100101011100100011;
        11'd1960: TDATA = 37'b0110001000101100110101001011100100001;
        11'd1961: TDATA = 37'b0110001001000011111101001011100100000;
        11'd1962: TDATA = 37'b0110001001011011000100101011100011110;
        11'd1963: TDATA = 37'b0110001001110010001100001011100011101;
        11'd1964: TDATA = 37'b0110001010001001010011001011100011011;
        11'd1965: TDATA = 37'b0110001010100000011001101011100011010;
        11'd1966: TDATA = 37'b0110001010110111100000001011100011000;
        11'd1967: TDATA = 37'b0110001011001110100101101011100010111;
        11'd1968: TDATA = 37'b0110001011100101101011001011100010101;
        11'd1969: TDATA = 37'b0110001011111100110000101011100010100;
        11'd1970: TDATA = 37'b0110001100010011110101001011100010010;
        11'd1971: TDATA = 37'b0110001100101010111001101011100010001;
        11'd1972: TDATA = 37'b0110001101000001111101101011100001111;
        11'd1973: TDATA = 37'b0110001101011001000001001011100001110;
        11'd1974: TDATA = 37'b0110001101110000000100001011100001100;
        11'd1975: TDATA = 37'b0110001110000111000111001011100001011;
        11'd1976: TDATA = 37'b0110001110011110001001101011100001001;
        11'd1977: TDATA = 37'b0110001110110101001011101011100001000;
        11'd1978: TDATA = 37'b0110001111001100001101101011100000110;
        11'd1979: TDATA = 37'b0110001111100011001111001011100000101;
        11'd1980: TDATA = 37'b0110001111111010010000001011100000011;
        11'd1981: TDATA = 37'b0110010000010001010000101011100000010;
        11'd1982: TDATA = 37'b0110010000101000010000101011100000000;
        11'd1983: TDATA = 37'b0110010000111111010000101011011111111;
        11'd1984: TDATA = 37'b0110010001010110010000001011011111101;
        11'd1985: TDATA = 37'b0110010001101101001111001011011111100;
        11'd1986: TDATA = 37'b0110010010000100001110001011011111010;
        11'd1987: TDATA = 37'b0110010010011011001100101011011111001;
        11'd1988: TDATA = 37'b0110010010110010001010101011011110111;
        11'd1989: TDATA = 37'b0110010011001001001000001011011110110;
        11'd1990: TDATA = 37'b0110010011100000000101101011011110100;
        11'd1991: TDATA = 37'b0110010011110111000010101011011110011;
        11'd1992: TDATA = 37'b0110010100001101111111001011011110001;
        11'd1993: TDATA = 37'b0110010100100100111011001011011110000;
        11'd1994: TDATA = 37'b0110010100111011110111001011011101111;
        11'd1995: TDATA = 37'b0110010101010010110010101011011101101;
        11'd1996: TDATA = 37'b0110010101101001101101101011011101100;
        11'd1997: TDATA = 37'b0110010110000000101000001011011101010;
        11'd1998: TDATA = 37'b0110010110010111100010101011011101001;
        11'd1999: TDATA = 37'b0110010110101110011100101011011100111;
        11'd2000: TDATA = 37'b0110010111000101010110001011011100110;
        11'd2001: TDATA = 37'b0110010111011100001111101011011100100;
        11'd2002: TDATA = 37'b0110010111110011001000001011011100011;
        11'd2003: TDATA = 37'b0110011000001010000000101011011100001;
        11'd2004: TDATA = 37'b0110011000100000111001001011011100000;
        11'd2005: TDATA = 37'b0110011000110111110000101011011011110;
        11'd2006: TDATA = 37'b0110011001001110101000001011011011101;
        11'd2007: TDATA = 37'b0110011001100101011111001011011011011;
        11'd2008: TDATA = 37'b0110011001111100010110001011011011010;
        11'd2009: TDATA = 37'b0110011010010011001100001011011011001;
        11'd2010: TDATA = 37'b0110011010101010000010001011011010111;
        11'd2011: TDATA = 37'b0110011011000000110111101011011010110;
        11'd2012: TDATA = 37'b0110011011010111101101001011011010100;
        11'd2013: TDATA = 37'b0110011011101110100010001011011010011;
        11'd2014: TDATA = 37'b0110011100000101010110101011011010001;
        11'd2015: TDATA = 37'b0110011100011100001010101011011010000;
        11'd2016: TDATA = 37'b0110011100110010111110001011011001110;
        11'd2017: TDATA = 37'b0110011101001001110001101011011001101;
        11'd2018: TDATA = 37'b0110011101100000100100101011011001100;
        11'd2019: TDATA = 37'b0110011101110111010111101011011001010;
        11'd2020: TDATA = 37'b0110011110001110001001101011011001001;
        11'd2021: TDATA = 37'b0110011110100100111011101011011000111;
        11'd2022: TDATA = 37'b0110011110111011101101101011011000110;
        11'd2023: TDATA = 37'b0110011111010010011110101011011000100;
        11'd2024: TDATA = 37'b0110011111101001001111101011011000011;
        11'd2025: TDATA = 37'b0110100000000000000000001011011000001;
        11'd2026: TDATA = 37'b0110100000010110110000001011011000000;
        11'd2027: TDATA = 37'b0110100000101101100000001011010111111;
        11'd2028: TDATA = 37'b0110100001000100001111101011010111101;
        11'd2029: TDATA = 37'b0110100001011010111110101011010111100;
        11'd2030: TDATA = 37'b0110100001110001101101101011010111010;
        11'd2031: TDATA = 37'b0110100010001000011011101011010111001;
        11'd2032: TDATA = 37'b0110100010011111001001101011010110111;
        11'd2033: TDATA = 37'b0110100010110101110111101011010110110;
        11'd2034: TDATA = 37'b0110100011001100100100101011010110101;
        11'd2035: TDATA = 37'b0110100011100011010001101011010110011;
        11'd2036: TDATA = 37'b0110100011111001111110001011010110010;
        11'd2037: TDATA = 37'b0110100100010000101010101011010110000;
        11'd2038: TDATA = 37'b0110100100100111010110101011010101111;
        11'd2039: TDATA = 37'b0110100100111110000010001011010101101;
        11'd2040: TDATA = 37'b0110100101010100101101001011010101100;
        11'd2041: TDATA = 37'b0110100101101011011000001011010101011;
        11'd2042: TDATA = 37'b0110100110000010000010101011010101001;
        11'd2043: TDATA = 37'b0110100110011000101100101011010101000;
        11'd2044: TDATA = 37'b0110100110101111010110001011010100110;
        11'd2045: TDATA = 37'b0110100111000101111111101011010100101;
        11'd2046: TDATA = 37'b0110100111011100101000101011010100011;
        11'd2047: TDATA = 37'b0110100111110011010001101011010100010;
        11'd0: TDATA = 37'b0110101000001001111001110110101000001;
        11'd1: TDATA = 37'b0110101000110111001001010110100111100;
        11'd2: TDATA = 37'b0110101001100100010111110110100110110;
        11'd3: TDATA = 37'b0110101010010001100100010110100110000;
        11'd4: TDATA = 37'b0110101010111110101111110110100101011;
        11'd5: TDATA = 37'b0110101011101011111001110110100100101;
        11'd6: TDATA = 37'b0110101100011001000010010110100011111;
        11'd7: TDATA = 37'b0110101101000110001001010110100011010;
        11'd8: TDATA = 37'b0110101101110011001111010110100010100;
        11'd9: TDATA = 37'b0110101110100000010011110110100001111;
        11'd10: TDATA = 37'b0110101111001101010110110110100001001;
        11'd11: TDATA = 37'b0110101111111010011000010110100000100;
        11'd12: TDATA = 37'b0110110000100111011000010110011111110;
        11'd13: TDATA = 37'b0110110001010100010111010110011111000;
        11'd14: TDATA = 37'b0110110010000001010100110110011110011;
        11'd15: TDATA = 37'b0110110010101110010000110110011101101;
        11'd16: TDATA = 37'b0110110011011011001011010110011101000;
        11'd17: TDATA = 37'b0110110100001000000100010110011100010;
        11'd18: TDATA = 37'b0110110100110100111100010110011011101;
        11'd19: TDATA = 37'b0110110101100001110010110110011010111;
        11'd20: TDATA = 37'b0110110110001110100111110110011010010;
        11'd21: TDATA = 37'b0110110110111011011011110110011001100;
        11'd22: TDATA = 37'b0110110111101000001110010110011000111;
        11'd23: TDATA = 37'b0110111000010100111111010110011000001;
        11'd24: TDATA = 37'b0110111001000001101110110110010111100;
        11'd25: TDATA = 37'b0110111001101110011100110110010110110;
        11'd26: TDATA = 37'b0110111010011011001001110110010110001;
        11'd27: TDATA = 37'b0110111011000111110101010110010101011;
        11'd28: TDATA = 37'b0110111011110100011111110110010100110;
        11'd29: TDATA = 37'b0110111100100001001000010110010100001;
        11'd30: TDATA = 37'b0110111101001101101111110110010011011;
        11'd31: TDATA = 37'b0110111101111010010110010110010010110;
        11'd32: TDATA = 37'b0110111110100110111010110110010010000;
        11'd33: TDATA = 37'b0110111111010011011110010110010001011;
        11'd34: TDATA = 37'b0111000000000000000000010110010000110;
        11'd35: TDATA = 37'b0111000000101100100000110110010000000;
        11'd36: TDATA = 37'b0111000001011001000000010110001111011;
        11'd37: TDATA = 37'b0111000010000101011110010110001110101;
        11'd38: TDATA = 37'b0111000010110001111011010110001110000;
        11'd39: TDATA = 37'b0111000011011110010110010110001101011;
        11'd40: TDATA = 37'b0111000100001010110000010110001100101;
        11'd41: TDATA = 37'b0111000100110111001001010110001100000;
        11'd42: TDATA = 37'b0111000101100011100000010110001011011;
        11'd43: TDATA = 37'b0111000110001111110110010110001010101;
        11'd44: TDATA = 37'b0111000110111100001011010110001010000;
        11'd45: TDATA = 37'b0111000111101000011110110110001001011;
        11'd46: TDATA = 37'b0111001000010100110000110110001000101;
        11'd47: TDATA = 37'b0111001001000001000001010110001000000;
        11'd48: TDATA = 37'b0111001001101101010000110110000111011;
        11'd49: TDATA = 37'b0111001010011001011110110110000110110;
        11'd50: TDATA = 37'b0111001011000101101011010110000110000;
        11'd51: TDATA = 37'b0111001011110001110110110110000101011;
        11'd52: TDATA = 37'b0111001100011110000000110110000100110;
        11'd53: TDATA = 37'b0111001101001010001001110110000100001;
        11'd54: TDATA = 37'b0111001101110110010001010110000011011;
        11'd55: TDATA = 37'b0111001110100010010111010110000010110;
        11'd56: TDATA = 37'b0111001111001110011100010110000010001;
        11'd57: TDATA = 37'b0111001111111010011111110110000001100;
        11'd58: TDATA = 37'b0111010000100110100010010110000000110;
        11'd59: TDATA = 37'b0111010001010010100011010110000000001;
        11'd60: TDATA = 37'b0111010001111110100010110101111111100;
        11'd61: TDATA = 37'b0111010010101010100001010101111110111;
        11'd62: TDATA = 37'b0111010011010110011110010101111110010;
        11'd63: TDATA = 37'b0111010100000010011001110101111101101;
        11'd64: TDATA = 37'b0111010100101110010100010101111100111;
        11'd65: TDATA = 37'b0111010101011010001101110101111100010;
        11'd66: TDATA = 37'b0111010110000110000101110101111011101;
        11'd67: TDATA = 37'b0111010110110001111100010101111011000;
        11'd68: TDATA = 37'b0111010111011101110001010101111010011;
        11'd69: TDATA = 37'b0111011000001001100101110101111001110;
        11'd70: TDATA = 37'b0111011000110101011000010101111001000;
        11'd71: TDATA = 37'b0111011001100001001001110101111000011;
        11'd72: TDATA = 37'b0111011010001100111001110101110111110;
        11'd73: TDATA = 37'b0111011010111000101000110101110111001;
        11'd74: TDATA = 37'b0111011011100100010110110101110110100;
        11'd75: TDATA = 37'b0111011100010000000010110101110101111;
        11'd76: TDATA = 37'b0111011100111011101101110101110101010;
        11'd77: TDATA = 37'b0111011101100111010111110101110100101;
        11'd78: TDATA = 37'b0111011110010011000000010101110100000;
        11'd79: TDATA = 37'b0111011110111110100111110101110011011;
        11'd80: TDATA = 37'b0111011111101010001101110101110010110;
        11'd81: TDATA = 37'b0111100000010101110010010101110010001;
        11'd82: TDATA = 37'b0111100001000001010101110101110001011;
        11'd83: TDATA = 37'b0111100001101100111000010101110000110;
        11'd84: TDATA = 37'b0111100010011000011001010101110000001;
        11'd85: TDATA = 37'b0111100011000011111000110101101111100;
        11'd86: TDATA = 37'b0111100011101111010111010101101110111;
        11'd87: TDATA = 37'b0111100100011010110100110101101110010;
        11'd88: TDATA = 37'b0111100101000110010000110101101101101;
        11'd89: TDATA = 37'b0111100101110001101011010101101101000;
        11'd90: TDATA = 37'b0111100110011101000100110101101100011;
        11'd91: TDATA = 37'b0111100111001000011101010101101011110;
        11'd92: TDATA = 37'b0111100111110011110100010101101011001;
        11'd93: TDATA = 37'b0111101000011111001001110101101010100;
        11'd94: TDATA = 37'b0111101001001010011110010101101010000;
        11'd95: TDATA = 37'b0111101001110101110001110101101001011;
        11'd96: TDATA = 37'b0111101010100001000011110101101000110;
        11'd97: TDATA = 37'b0111101011001100010100010101101000001;
        11'd98: TDATA = 37'b0111101011110111100011110101100111100;
        11'd99: TDATA = 37'b0111101100100010110010010101100110111;
        11'd100: TDATA = 37'b0111101101001101111111010101100110010;
        11'd101: TDATA = 37'b0111101101111001001011010101100101101;
        11'd102: TDATA = 37'b0111101110100100010101110101100101000;
        11'd103: TDATA = 37'b0111101111001111011111010101100100011;
        11'd104: TDATA = 37'b0111101111111010100111010101100011110;
        11'd105: TDATA = 37'b0111110000100101101110010101100011001;
        11'd106: TDATA = 37'b0111110001010000110011110101100010100;
        11'd107: TDATA = 37'b0111110001111011111000110101100010000;
        11'd108: TDATA = 37'b0111110010100110111011110101100001011;
        11'd109: TDATA = 37'b0111110011010001111101110101100000110;
        11'd110: TDATA = 37'b0111110011111100111110110101100000001;
        11'd111: TDATA = 37'b0111110100100111111110010101011111100;
        11'd112: TDATA = 37'b0111110101010010111100110101011110111;
        11'd113: TDATA = 37'b0111110101111101111010010101011110010;
        11'd114: TDATA = 37'b0111110110101000110110010101011101110;
        11'd115: TDATA = 37'b0111110111010011110000110101011101001;
        11'd116: TDATA = 37'b0111110111111110101010010101011100100;
        11'd117: TDATA = 37'b0111111000101001100010110101011011111;
        11'd118: TDATA = 37'b0111111001010100011010010101011011010;
        11'd119: TDATA = 37'b0111111001111111010000010101011010110;
        11'd120: TDATA = 37'b0111111010101010000100110101011010001;
        11'd121: TDATA = 37'b0111111011010100111000010101011001100;
        11'd122: TDATA = 37'b0111111011111111101010110101011000111;
        11'd123: TDATA = 37'b0111111100101010011100010101011000010;
        11'd124: TDATA = 37'b0111111101010101001100010101010111110;
        11'd125: TDATA = 37'b0111111101111111111010110101010111001;
        11'd126: TDATA = 37'b0111111110101010101000110101010110100;
        11'd127: TDATA = 37'b0111111111010101010100110101010101111;
        11'd128: TDATA = 37'b1000000000000000000000010101010101011;
        11'd129: TDATA = 37'b1000000000101010101010010101010100110;
        11'd130: TDATA = 37'b1000000001010101010011010101010100001;
        11'd131: TDATA = 37'b1000000001111111111010110101010011100;
        11'd132: TDATA = 37'b1000000010101010100001010101010011000;
        11'd133: TDATA = 37'b1000000011010101000110110101010010011;
        11'd134: TDATA = 37'b1000000011111111101010110101010001110;
        11'd135: TDATA = 37'b1000000100101010001101110101010001010;
        11'd136: TDATA = 37'b1000000101010100101111110101010000101;
        11'd137: TDATA = 37'b1000000101111111010000010101010000000;
        11'd138: TDATA = 37'b1000000110101001101111110101001111100;
        11'd139: TDATA = 37'b1000000111010100001110010101001110111;
        11'd140: TDATA = 37'b1000000111111110101011010101001110010;
        11'd141: TDATA = 37'b1000001000101001000111010101001101110;
        11'd142: TDATA = 37'b1000001001010011100010010101001101001;
        11'd143: TDATA = 37'b1000001001111101111011110101001100100;
        11'd144: TDATA = 37'b1000001010101000010100010101001100000;
        11'd145: TDATA = 37'b1000001011010010101011110101001011011;
        11'd146: TDATA = 37'b1000001011111101000001110101001010110;
        11'd147: TDATA = 37'b1000001100100111010110110101001010010;
        11'd148: TDATA = 37'b1000001101010001101010110101001001101;
        11'd149: TDATA = 37'b1000001101111011111101010101001001000;
        11'd150: TDATA = 37'b1000001110100110001110110101001000100;
        11'd151: TDATA = 37'b1000001111010000011111010101000111111;
        11'd152: TDATA = 37'b1000001111111010101110010101000111011;
        11'd153: TDATA = 37'b1000010000100100111100110101000110110;
        11'd154: TDATA = 37'b1000010001001111001001010101000110001;
        11'd155: TDATA = 37'b1000010001111001010101010101000101101;
        11'd156: TDATA = 37'b1000010010100011011111110101000101000;
        11'd157: TDATA = 37'b1000010011001101101001010101000100100;
        11'd158: TDATA = 37'b1000010011110111110001110101000011111;
        11'd159: TDATA = 37'b1000010100100001111000110101000011011;
        11'd160: TDATA = 37'b1000010101001011111111010101000010110;
        11'd161: TDATA = 37'b1000010101110110000011110101000010010;
        11'd162: TDATA = 37'b1000010110100000000111110101000001101;
        11'd163: TDATA = 37'b1000010111001010001010010101000001000;
        11'd164: TDATA = 37'b1000010111110100001100010101000000100;
        11'd165: TDATA = 37'b1000011000011110001100010100111111111;
        11'd166: TDATA = 37'b1000011001001000001011110100111111011;
        11'd167: TDATA = 37'b1000011001110010001001110100111110110;
        11'd168: TDATA = 37'b1000011010011100000110110100111110010;
        11'd169: TDATA = 37'b1000011011000110000010110100111101101;
        11'd170: TDATA = 37'b1000011011101111111101110100111101001;
        11'd171: TDATA = 37'b1000011100011001110111010100111100100;
        11'd172: TDATA = 37'b1000011101000011101111110100111100000;
        11'd173: TDATA = 37'b1000011101101101100111010100111011011;
        11'd174: TDATA = 37'b1000011110010111011101010100111010111;
        11'd175: TDATA = 37'b1000011111000001010010110100111010010;
        11'd176: TDATA = 37'b1000011111101011000110110100111001110;
        11'd177: TDATA = 37'b1000100000010100111001110100111001010;
        11'd178: TDATA = 37'b1000100000111110101011010100111000101;
        11'd179: TDATA = 37'b1000100001101000011100010100111000001;
        11'd180: TDATA = 37'b1000100010010010001011110100110111100;
        11'd181: TDATA = 37'b1000100010111011111010010100110111000;
        11'd182: TDATA = 37'b1000100011100101100111110100110110011;
        11'd183: TDATA = 37'b1000100100001111010011110100110101111;
        11'd184: TDATA = 37'b1000100100111000111111010100110101010;
        11'd185: TDATA = 37'b1000100101100010101001010100110100110;
        11'd186: TDATA = 37'b1000100110001100010010010100110100010;
        11'd187: TDATA = 37'b1000100110110101111001110100110011101;
        11'd188: TDATA = 37'b1000100111011111100000110100110011001;
        11'd189: TDATA = 37'b1000101000001001000110010100110010100;
        11'd190: TDATA = 37'b1000101000110010101010110100110010000;
        11'd191: TDATA = 37'b1000101001011100001110010100110001100;
        11'd192: TDATA = 37'b1000101010000101110000110100110000111;
        11'd193: TDATA = 37'b1000101010101111010010010100110000011;
        11'd194: TDATA = 37'b1000101011011000110010010100101111111;
        11'd195: TDATA = 37'b1000101100000010010001010100101111010;
        11'd196: TDATA = 37'b1000101100101011101111010100101110110;
        11'd197: TDATA = 37'b1000101101010101001100010100101110010;
        11'd198: TDATA = 37'b1000101101111110101000010100101101101;
        11'd199: TDATA = 37'b1000101110101000000010110100101101001;
        11'd200: TDATA = 37'b1000101111010001011100110100101100101;
        11'd201: TDATA = 37'b1000101111111010110101010100101100000;
        11'd202: TDATA = 37'b1000110000100100001100110100101011100;
        11'd203: TDATA = 37'b1000110001001101100011010100101011000;
        11'd204: TDATA = 37'b1000110001110110111000110100101010011;
        11'd205: TDATA = 37'b1000110010100000001100110100101001111;
        11'd206: TDATA = 37'b1000110011001001100000010100101001011;
        11'd207: TDATA = 37'b1000110011110010110010010100101000110;
        11'd208: TDATA = 37'b1000110100011100000011010100101000010;
        11'd209: TDATA = 37'b1000110101000101010011010100100111110;
        11'd210: TDATA = 37'b1000110101101110100010010100100111010;
        11'd211: TDATA = 37'b1000110110010111101111110100100110101;
        11'd212: TDATA = 37'b1000110111000000111100110100100110001;
        11'd213: TDATA = 37'b1000110111101010001000010100100101101;
        11'd214: TDATA = 37'b1000111000010011010011010100100101000;
        11'd215: TDATA = 37'b1000111000111100011100110100100100100;
        11'd216: TDATA = 37'b1000111001100101100101010100100100000;
        11'd217: TDATA = 37'b1000111010001110101100110100100011100;
        11'd218: TDATA = 37'b1000111010110111110011010100100010111;
        11'd219: TDATA = 37'b1000111011100000111000010100100010011;
        11'd220: TDATA = 37'b1000111100001001111100110100100001111;
        11'd221: TDATA = 37'b1000111100110010111111110100100001011;
        11'd222: TDATA = 37'b1000111101011100000010010100100000111;
        11'd223: TDATA = 37'b1000111110000101000011010100100000010;
        11'd224: TDATA = 37'b1000111110101110000011010100011111110;
        11'd225: TDATA = 37'b1000111111010111000010010100011111010;
        11'd226: TDATA = 37'b1001000000000000000000010100011110110;
        11'd227: TDATA = 37'b1001000000101000111101010100011110010;
        11'd228: TDATA = 37'b1001000001010001111001010100011101101;
        11'd229: TDATA = 37'b1001000001111010110011110100011101001;
        11'd230: TDATA = 37'b1001000010100011101101110100011100101;
        11'd231: TDATA = 37'b1001000011001100100110010100011100001;
        11'd232: TDATA = 37'b1001000011110101011110010100011011101;
        11'd233: TDATA = 37'b1001000100011110010100110100011011001;
        11'd234: TDATA = 37'b1001000101000111001010010100011010100;
        11'd235: TDATA = 37'b1001000101101111111110110100011010000;
        11'd236: TDATA = 37'b1001000110011000110010010100011001100;
        11'd237: TDATA = 37'b1001000111000001100100110100011001000;
        11'd238: TDATA = 37'b1001000111101010010110010100011000100;
        11'd239: TDATA = 37'b1001001000010011000110110100011000000;
        11'd240: TDATA = 37'b1001001000111011110110010100010111100;
        11'd241: TDATA = 37'b1001001001100100100100110100010110111;
        11'd242: TDATA = 37'b1001001010001101010001110100010110011;
        11'd243: TDATA = 37'b1001001010110101111110010100010101111;
        11'd244: TDATA = 37'b1001001011011110101001110100010101011;
        11'd245: TDATA = 37'b1001001100000111010011110100010100111;
        11'd246: TDATA = 37'b1001001100101111111100110100010100011;
        11'd247: TDATA = 37'b1001001101011000100101010100010011111;
        11'd248: TDATA = 37'b1001001110000001001100010100010011011;
        11'd249: TDATA = 37'b1001001110101001110010110100010010111;
        11'd250: TDATA = 37'b1001001111010010010111110100010010011;
        11'd251: TDATA = 37'b1001001111111010111011110100010001110;
        11'd252: TDATA = 37'b1001010000100011011110110100010001010;
        11'd253: TDATA = 37'b1001010001001100000000110100010000110;
        11'd254: TDATA = 37'b1001010001110100100010010100010000010;
        11'd255: TDATA = 37'b1001010010011101000010010100001111110;
        11'd256: TDATA = 37'b1001010011000101100001010100001111010;
        11'd257: TDATA = 37'b1001010011101101111111010100001110110;
        11'd258: TDATA = 37'b1001010100010110011100010100001110010;
        11'd259: TDATA = 37'b1001010100111110111000010100001101110;
        11'd260: TDATA = 37'b1001010101100111010011010100001101010;
        11'd261: TDATA = 37'b1001010110001111101101010100001100110;
        11'd262: TDATA = 37'b1001010110111000000110010100001100010;
        11'd263: TDATA = 37'b1001010111100000011110010100001011110;
        11'd264: TDATA = 37'b1001011000001000110101010100001011010;
        11'd265: TDATA = 37'b1001011000110001001011010100001010110;
        11'd266: TDATA = 37'b1001011001011001100000010100001010010;
        11'd267: TDATA = 37'b1001011010000001110100010100001001110;
        11'd268: TDATA = 37'b1001011010101010000111010100001001010;
        11'd269: TDATA = 37'b1001011011010010011001010100001000110;
        11'd270: TDATA = 37'b1001011011111010101010010100001000010;
        11'd271: TDATA = 37'b1001011100100010111010010100000111110;
        11'd272: TDATA = 37'b1001011101001011001001010100000111010;
        11'd273: TDATA = 37'b1001011101110011010111010100000110110;
        11'd274: TDATA = 37'b1001011110011011100100010100000110010;
        11'd275: TDATA = 37'b1001011111000011110000010100000101110;
        11'd276: TDATA = 37'b1001011111101011111011010100000101010;
        11'd277: TDATA = 37'b1001100000010100000101010100000100110;
        11'd278: TDATA = 37'b1001100000111100001110010100000100010;
        11'd279: TDATA = 37'b1001100001100100010110010100000011110;
        11'd280: TDATA = 37'b1001100010001100011101010100000011010;
        11'd281: TDATA = 37'b1001100010110100100011010100000010110;
        11'd282: TDATA = 37'b1001100011011100101000110100000010010;
        11'd283: TDATA = 37'b1001100100000100101100110100000001111;
        11'd284: TDATA = 37'b1001100100101100101111110100000001011;
        11'd285: TDATA = 37'b1001100101010100110010010100000000111;
        11'd286: TDATA = 37'b1001100101111100110011010100000000011;
        11'd287: TDATA = 37'b1001100110100100110011010011111111111;
        11'd288: TDATA = 37'b1001100111001100110010110011111111011;
        11'd289: TDATA = 37'b1001100111110100110000110011111110111;
        11'd290: TDATA = 37'b1001101000011100101110010011111110011;
        11'd291: TDATA = 37'b1001101001000100101010110011111101111;
        11'd292: TDATA = 37'b1001101001101100100101110011111101011;
        11'd293: TDATA = 37'b1001101010010100100000010011111101000;
        11'd294: TDATA = 37'b1001101010111100011001110011111100100;
        11'd295: TDATA = 37'b1001101011100100010010010011111100000;
        11'd296: TDATA = 37'b1001101100001100001001110011111011100;
        11'd297: TDATA = 37'b1001101100110100000000010011111011000;
        11'd298: TDATA = 37'b1001101101011011110101110011111010100;
        11'd299: TDATA = 37'b1001101110000011101010010011111010000;
        11'd300: TDATA = 37'b1001101110101011011101110011111001101;
        11'd301: TDATA = 37'b1001101111010011010000010011111001001;
        11'd302: TDATA = 37'b1001101111111011000010010011111000101;
        11'd303: TDATA = 37'b1001110000100010110010110011111000001;
        11'd304: TDATA = 37'b1001110001001010100010110011110111101;
        11'd305: TDATA = 37'b1001110001110010010001010011110111001;
        11'd306: TDATA = 37'b1001110010011001111111010011110110110;
        11'd307: TDATA = 37'b1001110011000001101100010011110110010;
        11'd308: TDATA = 37'b1001110011101001011000010011110101110;
        11'd309: TDATA = 37'b1001110100010001000011010011110101010;
        11'd310: TDATA = 37'b1001110100111000101101010011110100110;
        11'd311: TDATA = 37'b1001110101100000010110010011110100010;
        11'd312: TDATA = 37'b1001110110000111111110010011110011111;
        11'd313: TDATA = 37'b1001110110101111100101110011110011011;
        11'd314: TDATA = 37'b1001110111010111001011110011110010111;
        11'd315: TDATA = 37'b1001110111111110110001010011110010011;
        11'd316: TDATA = 37'b1001111000100110010101010011110010000;
        11'd317: TDATA = 37'b1001111001001101111000110011110001100;
        11'd318: TDATA = 37'b1001111001110101011011010011110001000;
        11'd319: TDATA = 37'b1001111010011100111100110011110000100;
        11'd320: TDATA = 37'b1001111011000100011101010011110000000;
        11'd321: TDATA = 37'b1001111011101011111101010011101111101;
        11'd322: TDATA = 37'b1001111100010011011011110011101111001;
        11'd323: TDATA = 37'b1001111100111010111001010011101110101;
        11'd324: TDATA = 37'b1001111101100010010110010011101110001;
        11'd325: TDATA = 37'b1001111110001001110010010011101101110;
        11'd326: TDATA = 37'b1001111110110001001101010011101101010;
        11'd327: TDATA = 37'b1001111111011000100111010011101100110;
        11'd328: TDATA = 37'b1010000000000000000000010011101100010;
        11'd329: TDATA = 37'b1010000000100111011000010011101011111;
        11'd330: TDATA = 37'b1010000001001110101111110011101011011;
        11'd331: TDATA = 37'b1010000001110110000101110011101010111;
        11'd332: TDATA = 37'b1010000010011101011011010011101010100;
        11'd333: TDATA = 37'b1010000011000100101111110011101010000;
        11'd334: TDATA = 37'b1010000011101100000011010011101001100;
        11'd335: TDATA = 37'b1010000100010011010101110011101001000;
        11'd336: TDATA = 37'b1010000100111010100111010011101000101;
        11'd337: TDATA = 37'b1010000101100001111000010011101000001;
        11'd338: TDATA = 37'b1010000110001001000111110011100111101;
        11'd339: TDATA = 37'b1010000110110000010110110011100111010;
        11'd340: TDATA = 37'b1010000111010111100100110011100110110;
        11'd341: TDATA = 37'b1010000111111110110001110011100110010;
        11'd342: TDATA = 37'b1010001000100101111101110011100101111;
        11'd343: TDATA = 37'b1010001001001101001001010011100101011;
        11'd344: TDATA = 37'b1010001001110100010011010011100100111;
        11'd345: TDATA = 37'b1010001010011011011100110011100100100;
        11'd346: TDATA = 37'b1010001011000010100101010011100100000;
        11'd347: TDATA = 37'b1010001011101001101100110011100011100;
        11'd348: TDATA = 37'b1010001100010000110011010011100011001;
        11'd349: TDATA = 37'b1010001100110111111001010011100010101;
        11'd350: TDATA = 37'b1010001101011110111110010011100010001;
        11'd351: TDATA = 37'b1010001110000110000001110011100001110;
        11'd352: TDATA = 37'b1010001110101101000100110011100001010;
        11'd353: TDATA = 37'b1010001111010100000110110011100000111;
        11'd354: TDATA = 37'b1010001111111011001000010011100000011;
        11'd355: TDATA = 37'b1010010000100010001000010011011111111;
        11'd356: TDATA = 37'b1010010001001001000111110011011111100;
        11'd357: TDATA = 37'b1010010001110000000110010011011111000;
        11'd358: TDATA = 37'b1010010010010111000011110011011110100;
        11'd359: TDATA = 37'b1010010010111110000000010011011110001;
        11'd360: TDATA = 37'b1010010011100100111100010011011101101;
        11'd361: TDATA = 37'b1010010100001011110111010011011101010;
        11'd362: TDATA = 37'b1010010100110010110001010011011100110;
        11'd363: TDATA = 37'b1010010101011001101010010011011100010;
        11'd364: TDATA = 37'b1010010110000000100010010011011011111;
        11'd365: TDATA = 37'b1010010110100111011001110011011011011;
        11'd366: TDATA = 37'b1010010111001110001111110011011011000;
        11'd367: TDATA = 37'b1010010111110101000101010011011010100;
        11'd368: TDATA = 37'b1010011000011011111001110011011010001;
        11'd369: TDATA = 37'b1010011001000010101101110011011001101;
        11'd370: TDATA = 37'b1010011001101001100000010011011001001;
        11'd371: TDATA = 37'b1010011010010000010010010011011000110;
        11'd372: TDATA = 37'b1010011010110111000011010011011000010;
        11'd373: TDATA = 37'b1010011011011101110011010011010111111;
        11'd374: TDATA = 37'b1010011100000100100010110011010111011;
        11'd375: TDATA = 37'b1010011100101011010001010011010111000;
        11'd376: TDATA = 37'b1010011101010001111110110011010110100;
        11'd377: TDATA = 37'b1010011101111000101011010011010110001;
        11'd378: TDATA = 37'b1010011110011111010110110011010101101;
        11'd379: TDATA = 37'b1010011111000110000001110011010101010;
        11'd380: TDATA = 37'b1010011111101100101011110011010100110;
        11'd381: TDATA = 37'b1010100000010011010100110011010100010;
        11'd382: TDATA = 37'b1010100000111001111100110011010011111;
        11'd383: TDATA = 37'b1010100001100000100100010011010011011;
        11'd384: TDATA = 37'b1010100010000111001010110011010011000;
        11'd385: TDATA = 37'b1010100010101101110000010011010010100;
        11'd386: TDATA = 37'b1010100011010100010100110011010010001;
        11'd387: TDATA = 37'b1010100011111010111000110011010001101;
        11'd388: TDATA = 37'b1010100100100001011011010011010001010;
        11'd389: TDATA = 37'b1010100101000111111101110011010000110;
        11'd390: TDATA = 37'b1010100101101110011110110011010000011;
        11'd391: TDATA = 37'b1010100110010100111110110011001111111;
        11'd392: TDATA = 37'b1010100110111011011110010011001111100;
        11'd393: TDATA = 37'b1010100111100001111100110011001111000;
        11'd394: TDATA = 37'b1010101000001000011010110011001110101;
        11'd395: TDATA = 37'b1010101000101110110111010011001110010;
        11'd396: TDATA = 37'b1010101001010101010011010011001101110;
        11'd397: TDATA = 37'b1010101001111011101110110011001101011;
        11'd398: TDATA = 37'b1010101010100010001000110011001100111;
        11'd399: TDATA = 37'b1010101011001000100010010011001100100;
        11'd400: TDATA = 37'b1010101011101110111010110011001100000;
        11'd401: TDATA = 37'b1010101100010101010010010011001011101;
        11'd402: TDATA = 37'b1010101100111011101001010011001011001;
        11'd403: TDATA = 37'b1010101101100001111110110011001010110;
        11'd404: TDATA = 37'b1010101110001000010011110011001010010;
        11'd405: TDATA = 37'b1010101110101110101000010011001001111;
        11'd406: TDATA = 37'b1010101111010100111011110011001001100;
        11'd407: TDATA = 37'b1010101111111011001110010011001001000;
        11'd408: TDATA = 37'b1010110000100001011111110011001000101;
        11'd409: TDATA = 37'b1010110001000111110000010011001000001;
        11'd410: TDATA = 37'b1010110001101110000000010011000111110;
        11'd411: TDATA = 37'b1010110010010100001111010011000111011;
        11'd412: TDATA = 37'b1010110010111010011101110011000110111;
        11'd413: TDATA = 37'b1010110011100000101010110011000110100;
        11'd414: TDATA = 37'b1010110100000110110111010011000110000;
        11'd415: TDATA = 37'b1010110100101101000011010011000101101;
        11'd416: TDATA = 37'b1010110101010011001101110011000101010;
        11'd417: TDATA = 37'b1010110101111001010111110011000100110;
        11'd418: TDATA = 37'b1010110110011111100000110011000100011;
        11'd419: TDATA = 37'b1010110111000101101001010011000011111;
        11'd420: TDATA = 37'b1010110111101011110000110011000011100;
        11'd421: TDATA = 37'b1010111000010001110111010011000011001;
        11'd422: TDATA = 37'b1010111000110111111100110011000010101;
        11'd423: TDATA = 37'b1010111001011110000001110011000010010;
        11'd424: TDATA = 37'b1010111010000100000101110011000001111;
        11'd425: TDATA = 37'b1010111010101010001001010011000001011;
        11'd426: TDATA = 37'b1010111011010000001011010011000001000;
        11'd427: TDATA = 37'b1010111011110110001100110011000000100;
        11'd428: TDATA = 37'b1010111100011100001101110011000000001;
        11'd429: TDATA = 37'b1010111101000010001101110010111111110;
        11'd430: TDATA = 37'b1010111101101000001100110010111111010;
        11'd431: TDATA = 37'b1010111110001110001010110010111110111;
        11'd432: TDATA = 37'b1010111110110100001000010010111110100;
        11'd433: TDATA = 37'b1010111111011010000100110010111110000;
        11'd434: TDATA = 37'b1011000000000000000000010010111101101;
        11'd435: TDATA = 37'b1011000000100101111011010010111101010;
        11'd436: TDATA = 37'b1011000001001011110101010010111100110;
        11'd437: TDATA = 37'b1011000001110001101110010010111100011;
        11'd438: TDATA = 37'b1011000010010111100110110010111100000;
        11'd439: TDATA = 37'b1011000010111101011110010010111011100;
        11'd440: TDATA = 37'b1011000011100011010100110010111011001;
        11'd441: TDATA = 37'b1011000100001001001010110010111010110;
        11'd442: TDATA = 37'b1011000100101110111111110010111010011;
        11'd443: TDATA = 37'b1011000101010100110011110010111001111;
        11'd444: TDATA = 37'b1011000101111010100111010010111001100;
        11'd445: TDATA = 37'b1011000110100000011001110010111001001;
        11'd446: TDATA = 37'b1011000111000110001011110010111000101;
        11'd447: TDATA = 37'b1011000111101011111100110010111000010;
        11'd448: TDATA = 37'b1011001000010001101100110010110111111;
        11'd449: TDATA = 37'b1011001000110111011011110010110111011;
        11'd450: TDATA = 37'b1011001001011101001010010010110111000;
        11'd451: TDATA = 37'b1011001010000010111000010010110110101;
        11'd452: TDATA = 37'b1011001010101000100100110010110110010;
        11'd453: TDATA = 37'b1011001011001110010000110010110101110;
        11'd454: TDATA = 37'b1011001011110011111100010010110101011;
        11'd455: TDATA = 37'b1011001100011001100110010010110101000;
        11'd456: TDATA = 37'b1011001100111111010000010010110100101;
        11'd457: TDATA = 37'b1011001101100100111000110010110100001;
        11'd458: TDATA = 37'b1011001110001010100000110010110011110;
        11'd459: TDATA = 37'b1011001110110000000111110010110011011;
        11'd460: TDATA = 37'b1011001111010101101110010010110011000;
        11'd461: TDATA = 37'b1011001111111011010011110010110010100;
        11'd462: TDATA = 37'b1011010000100000111000010010110010001;
        11'd463: TDATA = 37'b1011010001000110011100010010110001110;
        11'd464: TDATA = 37'b1011010001101011111111010010110001011;
        11'd465: TDATA = 37'b1011010010010001100001110010110000111;
        11'd466: TDATA = 37'b1011010010110111000010110010110000100;
        11'd467: TDATA = 37'b1011010011011100100011110010110000001;
        11'd468: TDATA = 37'b1011010100000010000011010010101111110;
        11'd469: TDATA = 37'b1011010100100111100010110010101111011;
        11'd470: TDATA = 37'b1011010101001101000000110010101110111;
        11'd471: TDATA = 37'b1011010101110010011110010010101110100;
        11'd472: TDATA = 37'b1011010110010111111010110010101110001;
        11'd473: TDATA = 37'b1011010110111101010110110010101101110;
        11'd474: TDATA = 37'b1011010111100010110001110010101101011;
        11'd475: TDATA = 37'b1011011000001000001011110010101100111;
        11'd476: TDATA = 37'b1011011000101101100101010010101100100;
        11'd477: TDATA = 37'b1011011001010010111101110010101100001;
        11'd478: TDATA = 37'b1011011001111000010101110010101011110;
        11'd479: TDATA = 37'b1011011010011101101100110010101011011;
        11'd480: TDATA = 37'b1011011011000011000011010010101010111;
        11'd481: TDATA = 37'b1011011011101000011000110010101010100;
        11'd482: TDATA = 37'b1011011100001101101101010010101010001;
        11'd483: TDATA = 37'b1011011100110011000001010010101001110;
        11'd484: TDATA = 37'b1011011101011000010100010010101001011;
        11'd485: TDATA = 37'b1011011101111101100110010010101001000;
        11'd486: TDATA = 37'b1011011110100010110111110010101000100;
        11'd487: TDATA = 37'b1011011111001000001000110010101000001;
        11'd488: TDATA = 37'b1011011111101101011000110010100111110;
        11'd489: TDATA = 37'b1011100000010010100111110010100111011;
        11'd490: TDATA = 37'b1011100000110111110110010010100111000;
        11'd491: TDATA = 37'b1011100001011101000011110010100110101;
        11'd492: TDATA = 37'b1011100010000010010000010010100110001;
        11'd493: TDATA = 37'b1011100010100111011100010010100101110;
        11'd494: TDATA = 37'b1011100011001100100111110010100101011;
        11'd495: TDATA = 37'b1011100011110001110001110010100101000;
        11'd496: TDATA = 37'b1011100100010110111011110010100100101;
        11'd497: TDATA = 37'b1011100100111100000100010010100100010;
        11'd498: TDATA = 37'b1011100101100001001100110010100011111;
        11'd499: TDATA = 37'b1011100110000110010011110010100011100;
        11'd500: TDATA = 37'b1011100110101011011010010010100011000;
        11'd501: TDATA = 37'b1011100111010000100000010010100010101;
        11'd502: TDATA = 37'b1011100111110101100100110010100010010;
        11'd503: TDATA = 37'b1011101000011010101001010010100001111;
        11'd504: TDATA = 37'b1011101000111111101100110010100001100;
        11'd505: TDATA = 37'b1011101001100100101111010010100001001;
        11'd506: TDATA = 37'b1011101010001001110001010010100000110;
        11'd507: TDATA = 37'b1011101010101110110010010010100000011;
        11'd508: TDATA = 37'b1011101011010011110010010010100000000;
        11'd509: TDATA = 37'b1011101011111000110001110010011111101;
        11'd510: TDATA = 37'b1011101100011101110000110010011111001;
        11'd511: TDATA = 37'b1011101101000010101110110010011110110;
        11'd512: TDATA = 37'b1011101101100111101011110010011110011;
        11'd513: TDATA = 37'b1011101110001100101000010010011110000;
        11'd514: TDATA = 37'b1011101110110001100011110010011101101;
        11'd515: TDATA = 37'b1011101111010110011110110010011101010;
        11'd516: TDATA = 37'b1011101111111011011001010010011100111;
        11'd517: TDATA = 37'b1011110000100000010010010010011100100;
        11'd518: TDATA = 37'b1011110001000101001011010010011100001;
        11'd519: TDATA = 37'b1011110001101010000010110010011011110;
        11'd520: TDATA = 37'b1011110010001110111001110010011011011;
        11'd521: TDATA = 37'b1011110010110011110000010010011011000;
        11'd522: TDATA = 37'b1011110011011000100101110010011010101;
        11'd523: TDATA = 37'b1011110011111101011010110010011010010;
        11'd524: TDATA = 37'b1011110100100010001110110010011001111;
        11'd525: TDATA = 37'b1011110101000111000001110010011001100;
        11'd526: TDATA = 37'b1011110101101011110100010010011001000;
        11'd527: TDATA = 37'b1011110110010000100110010010011000101;
        11'd528: TDATA = 37'b1011110110110101010111010010011000010;
        11'd529: TDATA = 37'b1011110111011010000111010010010111111;
        11'd530: TDATA = 37'b1011110111111110110110110010010111100;
        11'd531: TDATA = 37'b1011111000100011100101010010010111001;
        11'd532: TDATA = 37'b1011111001001000010011010010010110110;
        11'd533: TDATA = 37'b1011111001101101000000110010010110011;
        11'd534: TDATA = 37'b1011111010010001101101010010010110000;
        11'd535: TDATA = 37'b1011111010110110011000110010010101101;
        11'd536: TDATA = 37'b1011111011011011000011110010010101010;
        11'd537: TDATA = 37'b1011111011111111101101110010010100111;
        11'd538: TDATA = 37'b1011111100100100010111010010010100100;
        11'd539: TDATA = 37'b1011111101001001000000010010010100001;
        11'd540: TDATA = 37'b1011111101101101100111110010010011110;
        11'd541: TDATA = 37'b1011111110010010001111010010010011011;
        11'd542: TDATA = 37'b1011111110110110110101110010010011000;
        11'd543: TDATA = 37'b1011111111011011011011010010010010101;
        11'd544: TDATA = 37'b1100000000000000000000010010010010010;
        11'd545: TDATA = 37'b1100000000100100100100010010010001111;
        11'd546: TDATA = 37'b1100000001001001000111110010010001100;
        11'd547: TDATA = 37'b1100000001101101101010110010010001001;
        11'd548: TDATA = 37'b1100000010010010001100110010010000110;
        11'd549: TDATA = 37'b1100000010110110101101110010010000011;
        11'd550: TDATA = 37'b1100000011011011001110010010010000000;
        11'd551: TDATA = 37'b1100000011111111101110010010001111101;
        11'd552: TDATA = 37'b1100000100100100001100110010001111010;
        11'd553: TDATA = 37'b1100000101001000101011010010001111000;
        11'd554: TDATA = 37'b1100000101101101001000110010001110101;
        11'd555: TDATA = 37'b1100000110010001100101110010001110010;
        11'd556: TDATA = 37'b1100000110110110000001110010001101111;
        11'd557: TDATA = 37'b1100000111011010011100110010001101100;
        11'd558: TDATA = 37'b1100000111111110110111010010001101001;
        11'd559: TDATA = 37'b1100001000100011010001010010001100110;
        11'd560: TDATA = 37'b1100001001000111101010010010001100011;
        11'd561: TDATA = 37'b1100001001101100000010110010001100000;
        11'd562: TDATA = 37'b1100001010010000011010010010001011101;
        11'd563: TDATA = 37'b1100001010110100110001010010001011010;
        11'd564: TDATA = 37'b1100001011011001000111010010001010111;
        11'd565: TDATA = 37'b1100001011111101011100110010001010100;
        11'd566: TDATA = 37'b1100001100100001110001010010001010001;
        11'd567: TDATA = 37'b1100001101000110000101010010001001110;
        11'd568: TDATA = 37'b1100001101101010011000110010001001011;
        11'd569: TDATA = 37'b1100001110001110101011010010001001001;
        11'd570: TDATA = 37'b1100001110110010111100110010001000110;
        11'd571: TDATA = 37'b1100001111010111001101110010001000011;
        11'd572: TDATA = 37'b1100001111111011011110010010001000000;
        11'd573: TDATA = 37'b1100010000011111101101110010000111101;
        11'd574: TDATA = 37'b1100010001000011111100110010000111010;
        11'd575: TDATA = 37'b1100010001101000001010110010000110111;
        11'd576: TDATA = 37'b1100010010001100011000010010000110100;
        11'd577: TDATA = 37'b1100010010110000100100110010000110001;
        11'd578: TDATA = 37'b1100010011010100110000110010000101110;
        11'd579: TDATA = 37'b1100010011111000111100010010000101100;
        11'd580: TDATA = 37'b1100010100011101000110110010000101001;
        11'd581: TDATA = 37'b1100010101000001010000010010000100110;
        11'd582: TDATA = 37'b1100010101100101011001110010000100011;
        11'd583: TDATA = 37'b1100010110001001100001110010000100000;
        11'd584: TDATA = 37'b1100010110101101101001110010000011101;
        11'd585: TDATA = 37'b1100010111010001110000010010000011010;
        11'd586: TDATA = 37'b1100010111110101110110110010000010111;
        11'd587: TDATA = 37'b1100011000011001111100010010000010100;
        11'd588: TDATA = 37'b1100011000111110000000110010000010010;
        11'd589: TDATA = 37'b1100011001100010000100110010000001111;
        11'd590: TDATA = 37'b1100011010000110001000010010000001100;
        11'd591: TDATA = 37'b1100011010101010001010110010000001001;
        11'd592: TDATA = 37'b1100011011001110001100110010000000110;
        11'd593: TDATA = 37'b1100011011110010001101110010000000011;
        11'd594: TDATA = 37'b1100011100010110001110010010000000000;
        11'd595: TDATA = 37'b1100011100111010001110010001111111110;
        11'd596: TDATA = 37'b1100011101011110001101010001111111011;
        11'd597: TDATA = 37'b1100011110000010001011110001111111000;
        11'd598: TDATA = 37'b1100011110100110001001010001111110101;
        11'd599: TDATA = 37'b1100011111001010000110010001111110010;
        11'd600: TDATA = 37'b1100011111101110000010010001111101111;
        11'd601: TDATA = 37'b1100100000010001111101110001111101101;
        11'd602: TDATA = 37'b1100100000110101111000110001111101010;
        11'd603: TDATA = 37'b1100100001011001110010110001111100111;
        11'd604: TDATA = 37'b1100100001111101101100010001111100100;
        11'd605: TDATA = 37'b1100100010100001100100110001111100001;
        11'd606: TDATA = 37'b1100100011000101011100110001111011111;
        11'd607: TDATA = 37'b1100100011101001010100010001111011100;
        11'd608: TDATA = 37'b1100100100001101001010110001111011001;
        11'd609: TDATA = 37'b1100100100110001000000110001111010110;
        11'd610: TDATA = 37'b1100100101010100110101110001111010011;
        11'd611: TDATA = 37'b1100100101111000101010010001111010000;
        11'd612: TDATA = 37'b1100100110011100011101110001111001110;
        11'd613: TDATA = 37'b1100100111000000010001010001111001011;
        11'd614: TDATA = 37'b1100100111100100000011010001111001000;
        11'd615: TDATA = 37'b1100101000000111110101010001111000101;
        11'd616: TDATA = 37'b1100101000101011100110010001111000010;
        11'd617: TDATA = 37'b1100101001001111010110010001111000000;
        11'd618: TDATA = 37'b1100101001110011000101110001110111101;
        11'd619: TDATA = 37'b1100101010010110110100110001110111010;
        11'd620: TDATA = 37'b1100101010111010100010110001110110111;
        11'd621: TDATA = 37'b1100101011011110010000010001110110101;
        11'd622: TDATA = 37'b1100101100000001111101010001110110010;
        11'd623: TDATA = 37'b1100101100100101101001010001110101111;
        11'd624: TDATA = 37'b1100101101001001010100110001110101100;
        11'd625: TDATA = 37'b1100101101101100111111010001110101001;
        11'd626: TDATA = 37'b1100101110010000101001010001110100111;
        11'd627: TDATA = 37'b1100101110110100010010110001110100100;
        11'd628: TDATA = 37'b1100101111010111111011010001110100001;
        11'd629: TDATA = 37'b1100101111111011100011010001110011110;
        11'd630: TDATA = 37'b1100110000011111001010110001110011100;
        11'd631: TDATA = 37'b1100110001000010110001010001110011001;
        11'd632: TDATA = 37'b1100110001100110010111010001110010110;
        11'd633: TDATA = 37'b1100110010001001111100010001110010011;
        11'd634: TDATA = 37'b1100110010101101100000110001110010001;
        11'd635: TDATA = 37'b1100110011010001000100110001110001110;
        11'd636: TDATA = 37'b1100110011110100100111110001110001011;
        11'd637: TDATA = 37'b1100110100011000001010010001110001000;
        11'd638: TDATA = 37'b1100110100111011101011110001110000110;
        11'd639: TDATA = 37'b1100110101011111001100110001110000011;
        11'd640: TDATA = 37'b1100110110000010101101010001110000000;
        11'd641: TDATA = 37'b1100110110100110001101010001101111101;
        11'd642: TDATA = 37'b1100110111001001101100010001101111011;
        11'd643: TDATA = 37'b1100110111101101001010010001101111000;
        11'd644: TDATA = 37'b1100111000010000101000010001101110101;
        11'd645: TDATA = 37'b1100111000110100000101010001101110011;
        11'd646: TDATA = 37'b1100111001010111100001010001101110000;
        11'd647: TDATA = 37'b1100111001111010111100110001101101101;
        11'd648: TDATA = 37'b1100111010011110010111110001101101010;
        11'd649: TDATA = 37'b1100111011000001110010010001101101000;
        11'd650: TDATA = 37'b1100111011100101001011110001101100101;
        11'd651: TDATA = 37'b1100111100001000100100110001101100010;
        11'd652: TDATA = 37'b1100111100101011111100110001101100000;
        11'd653: TDATA = 37'b1100111101001111010100110001101011101;
        11'd654: TDATA = 37'b1100111101110010101011010001101011010;
        11'd655: TDATA = 37'b1100111110010110000001110001101011000;
        11'd656: TDATA = 37'b1100111110111001010111010001101010101;
        11'd657: TDATA = 37'b1100111111011100101100010001101010010;
        11'd658: TDATA = 37'b1101000000000000000000010001101001111;
        11'd659: TDATA = 37'b1101000000100011010011110001101001101;
        11'd660: TDATA = 37'b1101000001000110100110110001101001010;
        11'd661: TDATA = 37'b1101000001101001111000110001101000111;
        11'd662: TDATA = 37'b1101000010001101001010010001101000101;
        11'd663: TDATA = 37'b1101000010110000011011010001101000010;
        11'd664: TDATA = 37'b1101000011010011101011010001100111111;
        11'd665: TDATA = 37'b1101000011110110111010110001100111101;
        11'd666: TDATA = 37'b1101000100011010001001110001100111010;
        11'd667: TDATA = 37'b1101000100111101010111110001100110111;
        11'd668: TDATA = 37'b1101000101100000100101010001100110101;
        11'd669: TDATA = 37'b1101000110000011110010010001100110010;
        11'd670: TDATA = 37'b1101000110100110111110010001100101111;
        11'd671: TDATA = 37'b1101000111001010001001110001100101101;
        11'd672: TDATA = 37'b1101000111101101010100110001100101010;
        11'd673: TDATA = 37'b1101001000010000011110110001100100111;
        11'd674: TDATA = 37'b1101001000110011101000010001100100101;
        11'd675: TDATA = 37'b1101001001010110110001010001100100010;
        11'd676: TDATA = 37'b1101001001111001111001110001100011111;
        11'd677: TDATA = 37'b1101001010011101000001010001100011101;
        11'd678: TDATA = 37'b1101001011000000000111110001100011010;
        11'd679: TDATA = 37'b1101001011100011001110010001100011000;
        11'd680: TDATA = 37'b1101001100000110010011110001100010101;
        11'd681: TDATA = 37'b1101001100101001011000110001100010010;
        11'd682: TDATA = 37'b1101001101001100011100110001100010000;
        11'd683: TDATA = 37'b1101001101101111100000010001100001101;
        11'd684: TDATA = 37'b1101001110010010100011010001100001010;
        11'd685: TDATA = 37'b1101001110110101100101110001100001000;
        11'd686: TDATA = 37'b1101001111011000100111010001100000101;
        11'd687: TDATA = 37'b1101001111111011101000010001100000011;
        11'd688: TDATA = 37'b1101010000011110101000010001100000000;
        11'd689: TDATA = 37'b1101010001000001101000010001011111101;
        11'd690: TDATA = 37'b1101010001100100100111010001011111011;
        11'd691: TDATA = 37'b1101010010000111100101010001011111000;
        11'd692: TDATA = 37'b1101010010101010100011010001011110101;
        11'd693: TDATA = 37'b1101010011001101100000010001011110011;
        11'd694: TDATA = 37'b1101010011110000011100110001011110000;
        11'd695: TDATA = 37'b1101010100010011011000010001011101110;
        11'd696: TDATA = 37'b1101010100110110010011010001011101011;
        11'd697: TDATA = 37'b1101010101011001001101110001011101000;
        11'd698: TDATA = 37'b1101010101111100000111110001011100110;
        11'd699: TDATA = 37'b1101010110011111000000110001011100011;
        11'd700: TDATA = 37'b1101010111000001111001010001011100001;
        11'd701: TDATA = 37'b1101010111100100110001010001011011110;
        11'd702: TDATA = 37'b1101011000000111101000010001011011011;
        11'd703: TDATA = 37'b1101011000101010011110110001011011001;
        11'd704: TDATA = 37'b1101011001001101010100110001011010110;
        11'd705: TDATA = 37'b1101011001110000001001110001011010100;
        11'd706: TDATA = 37'b1101011010010010111110110001011010001;
        11'd707: TDATA = 37'b1101011010110101110010110001011001111;
        11'd708: TDATA = 37'b1101011011011000100101110001011001100;
        11'd709: TDATA = 37'b1101011011111011011000110001011001001;
        11'd710: TDATA = 37'b1101011100011110001010110001011000111;
        11'd711: TDATA = 37'b1101011101000000111100010001011000100;
        11'd712: TDATA = 37'b1101011101100011101100110001011000010;
        11'd713: TDATA = 37'b1101011110000110011100110001010111111;
        11'd714: TDATA = 37'b1101011110101001001100010001010111101;
        11'd715: TDATA = 37'b1101011111001011111011010001010111010;
        11'd716: TDATA = 37'b1101011111101110101001010001010111000;
        11'd717: TDATA = 37'b1101100000010001010110110001010110101;
        11'd718: TDATA = 37'b1101100000110100000011110001010110010;
        11'd719: TDATA = 37'b1101100001010110110000010001010110000;
        11'd720: TDATA = 37'b1101100001111001011011110001010101101;
        11'd721: TDATA = 37'b1101100010011100000110110001010101011;
        11'd722: TDATA = 37'b1101100010111110110001010001010101000;
        11'd723: TDATA = 37'b1101100011100001011010110001010100110;
        11'd724: TDATA = 37'b1101100100000100000100010001010100011;
        11'd725: TDATA = 37'b1101100100100110101100110001010100001;
        11'd726: TDATA = 37'b1101100101001001010100010001010011110;
        11'd727: TDATA = 37'b1101100101101011111011110001010011100;
        11'd728: TDATA = 37'b1101100110001110100010010001010011001;
        11'd729: TDATA = 37'b1101100110110001001000010001010010110;
        11'd730: TDATA = 37'b1101100111010011101101010001010010100;
        11'd731: TDATA = 37'b1101100111110110010010010001010010001;
        11'd732: TDATA = 37'b1101101000011000110110010001010001111;
        11'd733: TDATA = 37'b1101101000111011011001110001010001100;
        11'd734: TDATA = 37'b1101101001011101111100010001010001010;
        11'd735: TDATA = 37'b1101101010000000011110010001010000111;
        11'd736: TDATA = 37'b1101101010100010111111110001010000101;
        11'd737: TDATA = 37'b1101101011000101100000110001010000010;
        11'd738: TDATA = 37'b1101101011101000000001010001010000000;
        11'd739: TDATA = 37'b1101101100001010100000110001001111101;
        11'd740: TDATA = 37'b1101101100101100111111110001001111011;
        11'd741: TDATA = 37'b1101101101001111011110010001001111000;
        11'd742: TDATA = 37'b1101101101110001111100010001001110110;
        11'd743: TDATA = 37'b1101101110010100011001010001001110011;
        11'd744: TDATA = 37'b1101101110110110110101110001001110001;
        11'd745: TDATA = 37'b1101101111011001010001110001001101110;
        11'd746: TDATA = 37'b1101101111111011101100110001001101100;
        11'd747: TDATA = 37'b1101110000011110000111110001001101001;
        11'd748: TDATA = 37'b1101110001000000100001110001001100111;
        11'd749: TDATA = 37'b1101110001100010111010110001001100100;
        11'd750: TDATA = 37'b1101110010000101010011110001001100010;
        11'd751: TDATA = 37'b1101110010100111101011110001001011111;
        11'd752: TDATA = 37'b1101110011001010000011110001001011101;
        11'd753: TDATA = 37'b1101110011101100011010010001001011011;
        11'd754: TDATA = 37'b1101110100001110110000110001001011000;
        11'd755: TDATA = 37'b1101110100110001000110010001001010110;
        11'd756: TDATA = 37'b1101110101010011011011110001001010011;
        11'd757: TDATA = 37'b1101110101110101110000010001001010001;
        11'd758: TDATA = 37'b1101110110011000000011110001001001110;
        11'd759: TDATA = 37'b1101110110111010010111010001001001100;
        11'd760: TDATA = 37'b1101110111011100101001110001001001001;
        11'd761: TDATA = 37'b1101110111111110111011110001001000111;
        11'd762: TDATA = 37'b1101111000100001001101010001001000100;
        11'd763: TDATA = 37'b1101111001000011011101110001001000010;
        11'd764: TDATA = 37'b1101111001100101101110010001000111111;
        11'd765: TDATA = 37'b1101111010000111111101110001000111101;
        11'd766: TDATA = 37'b1101111010101010001100010001000111011;
        11'd767: TDATA = 37'b1101111011001100011010110001000111000;
        11'd768: TDATA = 37'b1101111011101110101000110001000110110;
        11'd769: TDATA = 37'b1101111100010000110101110001000110011;
        11'd770: TDATA = 37'b1101111100110011000010010001000110001;
        11'd771: TDATA = 37'b1101111101010101001101110001000101110;
        11'd772: TDATA = 37'b1101111101110111011001010001000101100;
        11'd773: TDATA = 37'b1101111110011001100011110001000101001;
        11'd774: TDATA = 37'b1101111110111011101101110001000100111;
        11'd775: TDATA = 37'b1101111111011101110111010001000100101;
        11'd776: TDATA = 37'b1110000000000000000000010001000100010;
        11'd777: TDATA = 37'b1110000000100010001000010001000100000;
        11'd778: TDATA = 37'b1110000001000100010000010001000011101;
        11'd779: TDATA = 37'b1110000001100110010111010001000011011;
        11'd780: TDATA = 37'b1110000010001000011101110001000011000;
        11'd781: TDATA = 37'b1110000010101010100011010001000010110;
        11'd782: TDATA = 37'b1110000011001100101000110001000010100;
        11'd783: TDATA = 37'b1110000011101110101101010001000010001;
        11'd784: TDATA = 37'b1110000100010000110001010001000001111;
        11'd785: TDATA = 37'b1110000100110010110100110001000001100;
        11'd786: TDATA = 37'b1110000101010100110111010001000001010;
        11'd787: TDATA = 37'b1110000101110110111001110001000001000;
        11'd788: TDATA = 37'b1110000110011000111011010001000000101;
        11'd789: TDATA = 37'b1110000110111010111100010001000000011;
        11'd790: TDATA = 37'b1110000111011100111100010001000000000;
        11'd791: TDATA = 37'b1110000111111110111100010000111111110;
        11'd792: TDATA = 37'b1110001000100000111011010000111111100;
        11'd793: TDATA = 37'b1110001001000010111010010000111111001;
        11'd794: TDATA = 37'b1110001001100100111000010000111110111;
        11'd795: TDATA = 37'b1110001010000110110101010000111110100;
        11'd796: TDATA = 37'b1110001010101000110010010000111110010;
        11'd797: TDATA = 37'b1110001011001010101110010000111110000;
        11'd798: TDATA = 37'b1110001011101100101010010000111101101;
        11'd799: TDATA = 37'b1110001100001110100101010000111101011;
        11'd800: TDATA = 37'b1110001100110000011111010000111101000;
        11'd801: TDATA = 37'b1110001101010010011001010000111100110;
        11'd802: TDATA = 37'b1110001101110100010010010000111100100;
        11'd803: TDATA = 37'b1110001110010110001011010000111100001;
        11'd804: TDATA = 37'b1110001110111000000011010000111011111;
        11'd805: TDATA = 37'b1110001111011001111010110000111011101;
        11'd806: TDATA = 37'b1110001111111011110001010000111011010;
        11'd807: TDATA = 37'b1110010000011101100111110000111011000;
        11'd808: TDATA = 37'b1110010000111111011101010000111010101;
        11'd809: TDATA = 37'b1110010001100001010010010000111010011;
        11'd810: TDATA = 37'b1110010010000011000110110000111010001;
        11'd811: TDATA = 37'b1110010010100100111010110000111001110;
        11'd812: TDATA = 37'b1110010011000110101110010000111001100;
        11'd813: TDATA = 37'b1110010011101000100000110000111001010;
        11'd814: TDATA = 37'b1110010100001010010010110000111000111;
        11'd815: TDATA = 37'b1110010100101100000100110000111000101;
        11'd816: TDATA = 37'b1110010101001101110101010000111000011;
        11'd817: TDATA = 37'b1110010101101111100101110000111000000;
        11'd818: TDATA = 37'b1110010110010001010101110000110111110;
        11'd819: TDATA = 37'b1110010110110011000100110000110111100;
        11'd820: TDATA = 37'b1110010111010100110011010000110111001;
        11'd821: TDATA = 37'b1110010111110110100001010000110110111;
        11'd822: TDATA = 37'b1110011000011000001110110000110110101;
        11'd823: TDATA = 37'b1110011000111001111011110000110110010;
        11'd824: TDATA = 37'b1110011001011011100111110000110110000;
        11'd825: TDATA = 37'b1110011001111101010011110000110101110;
        11'd826: TDATA = 37'b1110011010011110111110110000110101011;
        11'd827: TDATA = 37'b1110011011000000101001010000110101001;
        11'd828: TDATA = 37'b1110011011100010010011010000110100111;
        11'd829: TDATA = 37'b1110011100000011111100110000110100100;
        11'd830: TDATA = 37'b1110011100100101100101010000110100010;
        11'd831: TDATA = 37'b1110011101000111001101110000110100000;
        11'd832: TDATA = 37'b1110011101101000110101010000110011101;
        11'd833: TDATA = 37'b1110011110001010011100010000110011011;
        11'd834: TDATA = 37'b1110011110101100000010110000110011001;
        11'd835: TDATA = 37'b1110011111001101101000110000110010110;
        11'd836: TDATA = 37'b1110011111101111001101110000110010100;
        11'd837: TDATA = 37'b1110100000010000110010110000110010010;
        11'd838: TDATA = 37'b1110100000110010010110110000110001111;
        11'd839: TDATA = 37'b1110100001010011111010010000110001101;
        11'd840: TDATA = 37'b1110100001110101011101010000110001011;
        11'd841: TDATA = 37'b1110100010010110111111110000110001001;
        11'd842: TDATA = 37'b1110100010111000100001010000110000110;
        11'd843: TDATA = 37'b1110100011011010000010110000110000100;
        11'd844: TDATA = 37'b1110100011111011100011010000110000010;
        11'd845: TDATA = 37'b1110100100011101000011110000101111111;
        11'd846: TDATA = 37'b1110100100111110100011010000101111101;
        11'd847: TDATA = 37'b1110100101100000000010010000101111011;
        11'd848: TDATA = 37'b1110100110000001100000010000101111000;
        11'd849: TDATA = 37'b1110100110100010111110010000101110110;
        11'd850: TDATA = 37'b1110100111000100011011110000101110100;
        11'd851: TDATA = 37'b1110100111100101111000010000101110010;
        11'd852: TDATA = 37'b1110101000000111010100010000101101111;
        11'd853: TDATA = 37'b1110101000101000101111110000101101101;
        11'd854: TDATA = 37'b1110101001001010001010110000101101011;
        11'd855: TDATA = 37'b1110101001101011100101010000101101000;
        11'd856: TDATA = 37'b1110101010001100111111010000101100110;
        11'd857: TDATA = 37'b1110101010101110011000010000101100100;
        11'd858: TDATA = 37'b1110101011001111110001010000101100010;
        11'd859: TDATA = 37'b1110101011110001001001010000101011111;
        11'd860: TDATA = 37'b1110101100010010100000110000101011101;
        11'd861: TDATA = 37'b1110101100110011110111110000101011011;
        11'd862: TDATA = 37'b1110101101010101001110010000101011001;
        11'd863: TDATA = 37'b1110101101110110100100010000101010110;
        11'd864: TDATA = 37'b1110101110010111111001010000101010100;
        11'd865: TDATA = 37'b1110101110111001001110010000101010010;
        11'd866: TDATA = 37'b1110101111011010100010010000101010000;
        11'd867: TDATA = 37'b1110101111111011110101110000101001101;
        11'd868: TDATA = 37'b1110110000011101001000110000101001011;
        11'd869: TDATA = 37'b1110110000111110011011010000101001001;
        11'd870: TDATA = 37'b1110110001011111101101010000101000111;
        11'd871: TDATA = 37'b1110110010000000111110110000101000100;
        11'd872: TDATA = 37'b1110110010100010001111010000101000010;
        11'd873: TDATA = 37'b1110110011000011011111110000101000000;
        11'd874: TDATA = 37'b1110110011100100101111010000100111110;
        11'd875: TDATA = 37'b1110110100000101111110010000100111011;
        11'd876: TDATA = 37'b1110110100100111001100110000100111001;
        11'd877: TDATA = 37'b1110110101001000011010110000100110111;
        11'd878: TDATA = 37'b1110110101101001101000010000100110101;
        11'd879: TDATA = 37'b1110110110001010110101010000100110010;
        11'd880: TDATA = 37'b1110110110101100000001110000100110000;
        11'd881: TDATA = 37'b1110110111001101001101010000100101110;
        11'd882: TDATA = 37'b1110110111101110011000110000100101100;
        11'd883: TDATA = 37'b1110111000001111100011010000100101001;
        11'd884: TDATA = 37'b1110111000110000101101010000100100111;
        11'd885: TDATA = 37'b1110111001010001110110110000100100101;
        11'd886: TDATA = 37'b1110111001110010111111110000100100011;
        11'd887: TDATA = 37'b1110111010010100001000010000100100001;
        11'd888: TDATA = 37'b1110111010110101010000010000100011110;
        11'd889: TDATA = 37'b1110111011010110010111010000100011100;
        11'd890: TDATA = 37'b1110111011110111011110010000100011010;
        11'd891: TDATA = 37'b1110111100011000100100010000100011000;
        11'd892: TDATA = 37'b1110111100111001101001110000100010101;
        11'd893: TDATA = 37'b1110111101011010101111010000100010011;
        11'd894: TDATA = 37'b1110111101111011110011110000100010001;
        11'd895: TDATA = 37'b1110111110011100110111110000100001111;
        11'd896: TDATA = 37'b1110111110111101111011010000100001101;
        11'd897: TDATA = 37'b1110111111011110111101110000100001010;
        11'd898: TDATA = 37'b1111000000000000000000010000100001000;
        11'd899: TDATA = 37'b1111000000100001000010010000100000110;
        11'd900: TDATA = 37'b1111000001000010000011010000100000100;
        11'd901: TDATA = 37'b1111000001100011000011110000100000010;
        11'd902: TDATA = 37'b1111000010000100000100010000011111111;
        11'd903: TDATA = 37'b1111000010100101000011110000011111101;
        11'd904: TDATA = 37'b1111000011000110000010110000011111011;
        11'd905: TDATA = 37'b1111000011100111000001010000011111001;
        11'd906: TDATA = 37'b1111000100000111111111010000011110111;
        11'd907: TDATA = 37'b1111000100101000111100110000011110101;
        11'd908: TDATA = 37'b1111000101001001111001010000011110010;
        11'd909: TDATA = 37'b1111000101101010110101110000011110000;
        11'd910: TDATA = 37'b1111000110001011110001110000011101110;
        11'd911: TDATA = 37'b1111000110101100101100110000011101100;
        11'd912: TDATA = 37'b1111000111001101100111010000011101010;
        11'd913: TDATA = 37'b1111000111101110100001110000011100111;
        11'd914: TDATA = 37'b1111001000001111011011010000011100101;
        11'd915: TDATA = 37'b1111001000110000010100010000011100011;
        11'd916: TDATA = 37'b1111001001010001001100110000011100001;
        11'd917: TDATA = 37'b1111001001110010000100110000011011111;
        11'd918: TDATA = 37'b1111001010010010111100010000011011101;
        11'd919: TDATA = 37'b1111001010110011110010110000011011010;
        11'd920: TDATA = 37'b1111001011010100101001010000011011000;
        11'd921: TDATA = 37'b1111001011110101011111010000011010110;
        11'd922: TDATA = 37'b1111001100010110010100010000011010100;
        11'd923: TDATA = 37'b1111001100110111001001010000011010010;
        11'd924: TDATA = 37'b1111001101010111111101010000011010000;
        11'd925: TDATA = 37'b1111001101111000110000110000011001101;
        11'd926: TDATA = 37'b1111001110011001100100010000011001011;
        11'd927: TDATA = 37'b1111001110111010010110110000011001001;
        11'd928: TDATA = 37'b1111001111011011001000110000011000111;
        11'd929: TDATA = 37'b1111001111111011111010010000011000101;
        11'd930: TDATA = 37'b1111010000011100101011010000011000011;
        11'd931: TDATA = 37'b1111010000111101011011010000011000001;
        11'd932: TDATA = 37'b1111010001011110001011010000010111110;
        11'd933: TDATA = 37'b1111010001111110111010110000010111100;
        11'd934: TDATA = 37'b1111010010011111101001010000010111010;
        11'd935: TDATA = 37'b1111010011000000010111110000010111000;
        11'd936: TDATA = 37'b1111010011100001000101110000010110110;
        11'd937: TDATA = 37'b1111010100000001110010110000010110100;
        11'd938: TDATA = 37'b1111010100100010011111010000010110010;
        11'd939: TDATA = 37'b1111010101000011001011110000010101111;
        11'd940: TDATA = 37'b1111010101100011110111010000010101101;
        11'd941: TDATA = 37'b1111010110000100100010010000010101011;
        11'd942: TDATA = 37'b1111010110100101001100110000010101001;
        11'd943: TDATA = 37'b1111010111000101110110110000010100111;
        11'd944: TDATA = 37'b1111010111100110100000010000010100101;
        11'd945: TDATA = 37'b1111011000000111001001010000010100011;
        11'd946: TDATA = 37'b1111011000100111110001110000010100001;
        11'd947: TDATA = 37'b1111011001001000011001010000010011110;
        11'd948: TDATA = 37'b1111011001101001000000110000010011100;
        11'd949: TDATA = 37'b1111011010001001100111110000010011010;
        11'd950: TDATA = 37'b1111011010101010001101110000010011000;
        11'd951: TDATA = 37'b1111011011001010110011110000010010110;
        11'd952: TDATA = 37'b1111011011101011011000110000010010100;
        11'd953: TDATA = 37'b1111011100001011111101110000010010010;
        11'd954: TDATA = 37'b1111011100101100100001110000010010000;
        11'd955: TDATA = 37'b1111011101001101000101110000010001110;
        11'd956: TDATA = 37'b1111011101101101101000110000010001011;
        11'd957: TDATA = 37'b1111011110001110001011010000010001001;
        11'd958: TDATA = 37'b1111011110101110101101010000010000111;
        11'd959: TDATA = 37'b1111011111001111001110110000010000101;
        11'd960: TDATA = 37'b1111011111101111101111110000010000011;
        11'd961: TDATA = 37'b1111100000010000010000010000010000001;
        11'd962: TDATA = 37'b1111100000110000110000010000001111111;
        11'd963: TDATA = 37'b1111100001010001001111110000001111101;
        11'd964: TDATA = 37'b1111100001110001101110110000001111011;
        11'd965: TDATA = 37'b1111100010010010001101010000001111001;
        11'd966: TDATA = 37'b1111100010110010101011010000001110111;
        11'd967: TDATA = 37'b1111100011010011001000010000001110100;
        11'd968: TDATA = 37'b1111100011110011100101010000001110010;
        11'd969: TDATA = 37'b1111100100010100000001110000001110000;
        11'd970: TDATA = 37'b1111100100110100011101010000001101110;
        11'd971: TDATA = 37'b1111100101010100111000110000001101100;
        11'd972: TDATA = 37'b1111100101110101010011110000001101010;
        11'd973: TDATA = 37'b1111100110010101101101110000001101000;
        11'd974: TDATA = 37'b1111100110110110000111110000001100110;
        11'd975: TDATA = 37'b1111100111010110100000110000001100100;
        11'd976: TDATA = 37'b1111100111110110111001010000001100010;
        11'd977: TDATA = 37'b1111101000010111010001110000001100000;
        11'd978: TDATA = 37'b1111101000110111101001010000001011110;
        11'd979: TDATA = 37'b1111101001011000000000010000001011100;
        11'd980: TDATA = 37'b1111101001111000010110110000001011001;
        11'd981: TDATA = 37'b1111101010011000101101010000001010111;
        11'd982: TDATA = 37'b1111101010111001000010110000001010101;
        11'd983: TDATA = 37'b1111101011011001010111110000001010011;
        11'd984: TDATA = 37'b1111101011111001101100010000001010001;
        11'd985: TDATA = 37'b1111101100011010000000010000001001111;
        11'd986: TDATA = 37'b1111101100111010010011110000001001101;
        11'd987: TDATA = 37'b1111101101011010100110110000001001011;
        11'd988: TDATA = 37'b1111101101111010111001010000001001001;
        11'd989: TDATA = 37'b1111101110011011001011010000001000111;
        11'd990: TDATA = 37'b1111101110111011011100110000001000101;
        11'd991: TDATA = 37'b1111101111011011101101110000001000011;
        11'd992: TDATA = 37'b1111101111111011111110010000001000001;
        11'd993: TDATA = 37'b1111110000011100001110010000000111111;
        11'd994: TDATA = 37'b1111110000111100011101110000000111101;
        11'd995: TDATA = 37'b1111110001011100101100010000000111011;
        11'd996: TDATA = 37'b1111110001111100111010110000000111001;
        11'd997: TDATA = 37'b1111110010011101001000110000000110111;
        11'd998: TDATA = 37'b1111110010111101010110010000000110101;
        11'd999: TDATA = 37'b1111110011011101100011010000000110010;
        11'd1000: TDATA = 37'b1111110011111101101111010000000110000;
        11'd1001: TDATA = 37'b1111110100011101111011010000000101110;
        11'd1002: TDATA = 37'b1111110100111110000110110000000101100;
        11'd1003: TDATA = 37'b1111110101011110010001010000000101010;
        11'd1004: TDATA = 37'b1111110101111110011011110000000101000;
        11'd1005: TDATA = 37'b1111110110011110100101110000000100110;
        11'd1006: TDATA = 37'b1111110110111110101110110000000100100;
        11'd1007: TDATA = 37'b1111110111011110110111110000000100010;
        11'd1008: TDATA = 37'b1111110111111110111111110000000100000;
        11'd1009: TDATA = 37'b1111111000011111000111110000000011110;
        11'd1010: TDATA = 37'b1111111000111111001111010000000011100;
        11'd1011: TDATA = 37'b1111111001011111010101110000000011010;
        11'd1012: TDATA = 37'b1111111001111111011100010000000011000;
        11'd1013: TDATA = 37'b1111111010011111100001110000000010110;
        11'd1014: TDATA = 37'b1111111010111111100111010000000010100;
        11'd1015: TDATA = 37'b1111111011011111101011110000000010010;
        11'd1016: TDATA = 37'b1111111011111111110000010000000010000;
        11'd1017: TDATA = 37'b1111111100011111110011110000000001110;
        11'd1018: TDATA = 37'b1111111100111111110111010000000001100;
        11'd1019: TDATA = 37'b1111111101011111111001110000000001010;
        11'd1020: TDATA = 37'b1111111101111111111100010000000001000;
        11'd1021: TDATA = 37'b1111111110011111111101110000000000110;
        11'd1022: TDATA = 37'b1111111110111111111111010000000000100;
        11'd1023: TDATA = 37'b1111111111011111111111110000000000010;
        endcase
    end
    endfunction

    wire [7:0] ex;
    wire [22:0] mx;
    assign ex = x[30:23];
    assign mx = x[22:0];
    
    wire [10:0] key;
    wire [12:0] h;
    assign key = x[23:13];
    assign h = x[12:0];

    wire [36:0] tdata;
    assign tdata = TDATA(key);

    wire [22:0] rtx0;
    wire [13:0] rtx0_inv;
    assign rtx0 = tdata[36:14];
    assign rtx0_inv = tdata[13:0];

    wire [7:0] ey;
    assign ey = (ex == 0) ? 0: 8'd63 + ex[7:1] + ex[0];

    wire [36:0] my_extend;
    assign my_extend = {rtx0,14'b0} + rtx0_inv * h;

    wire [22:0] my;
    assign my = my_extend[36:14];

    assign y = {1'b0,ey,my};

endmodule

