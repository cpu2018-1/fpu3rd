module fsqrt(
    input wire [31:0] x,
    output wire [31:0] y,
    input wire clk,
    input wire rstn);

    function [38:0] TDATA (
	input [9:0] INDEX
    );
    begin
	casex(INDEX)
        10'd0: TDATA = 39'b100001111011010101101001100011000100001;
        10'd1: TDATA = 39'b100001111001000101101000011011001101000;
        10'd2: TDATA = 39'b100001110111001101100111011111011011110;
        10'd3: TDATA = 39'b100001110100111101100110010111110110001;
        10'd4: TDATA = 39'b100001110010101101100101010000011010001;
        10'd5: TDATA = 39'b100001110000110101100100010100111111010;
        10'd6: TDATA = 39'b100001101110100101100011001101110100101;
        10'd7: TDATA = 39'b100001101100101101100010010010101000010;
        10'd8: TDATA = 39'b100001101010011101100001001011101111000;
        10'd9: TDATA = 39'b100001101000100101100000010000110001001;
        10'd10: TDATA = 39'b100001100110010101011111001010001001010;
        10'd11: TDATA = 39'b100001100100011101011110001111011001111;
        10'd12: TDATA = 39'b100001100010001101011101001001000011010;
        10'd13: TDATA = 39'b100001100000010101011100001110100010010;
        10'd14: TDATA = 39'b100001011110000101011011001000011100111;
        10'd15: TDATA = 39'b100001011100001101011010001110001010011;
        10'd16: TDATA = 39'b100001011001111101011001001000010110010;
        10'd17: TDATA = 39'b100001011000000101011000001110010010000;
        10'd18: TDATA = 39'b100001010110001101010111010100010100010;
        10'd19: TDATA = 39'b100001010011111101010110001110111001010;
        10'd20: TDATA = 39'b100001010010000101010101010101001001111;
        10'd21: TDATA = 39'b100001010000001101010100011011100001000;
        10'd22: TDATA = 39'b100001001101111101010011010110011110111;
        10'd23: TDATA = 39'b100001001100000101010010011101000100010;
        10'd24: TDATA = 39'b100001001010001101010001100011110000001;
        10'd25: TDATA = 39'b100001001000010101010000101010100010100;
        10'd26: TDATA = 39'b100001000110000101001111100110000001000;
        10'd27: TDATA = 39'b100001000100001101001110101101000001101;
        10'd28: TDATA = 39'b100001000010010101001101110100001000101;
        10'd29: TDATA = 39'b100001000000011101001100111011010110001;
        10'd30: TDATA = 39'b100000111110001101001011110111010101010;
        10'd31: TDATA = 39'b100000111100010101001010111110110000111;
        10'd32: TDATA = 39'b100000111010011101001010000110010011000;
        10'd33: TDATA = 39'b100000111000100101001001001101111011100;
        10'd34: TDATA = 39'b100000110110101101001000010101101010100;
        10'd35: TDATA = 39'b100000110100110101000111011101011111110;
        10'd36: TDATA = 39'b100000110010111101000110100101011011101;
        10'd37: TDATA = 39'b100000110000101101000101100010010010001;
        10'd38: TDATA = 39'b100000101110110101000100101010011100000;
        10'd39: TDATA = 39'b100000101100111101000011110010101100010;
        10'd40: TDATA = 39'b100000101011000101000010111011000010111;
        10'd41: TDATA = 39'b100000101001001101000010000011011111111;
        10'd42: TDATA = 39'b100000100111010101000001001100000011011;
        10'd43: TDATA = 39'b100000100101011101000000010100101101001;
        10'd44: TDATA = 39'b100000100011100100111111011101011101010;
        10'd45: TDATA = 39'b100000100001101100111110100110010011110;
        10'd46: TDATA = 39'b100000011111110100111101101111010000100;
        10'd47: TDATA = 39'b100000011101111100111100111000010011110;
        10'd48: TDATA = 39'b100000011100000100111100000001011101010;
        10'd49: TDATA = 39'b100000011010001100111011001010101101001;
        10'd50: TDATA = 39'b100000011000010100111010010100000011010;
        10'd51: TDATA = 39'b100000010110110100111001101000011001101;
        10'd52: TDATA = 39'b100000010100111100111000110001111011001;
        10'd53: TDATA = 39'b100000010011000100110111111011100011001;
        10'd54: TDATA = 39'b100000010001001100110111000101010001010;
        10'd55: TDATA = 39'b100000001111010100110110001111000101110;
        10'd56: TDATA = 39'b100000001101011100110101011001000000100;
        10'd57: TDATA = 39'b100000001011100100110100100011000001101;
        10'd58: TDATA = 39'b100000001010000100110011110111111010010;
        10'd59: TDATA = 39'b100000001000001100110011000010000110101;
        10'd60: TDATA = 39'b100000000110010100110010001100011001010;
        10'd61: TDATA = 39'b100000000100011100110001010110110010010;
        10'd62: TDATA = 39'b100000000010100100110000100001010001011;
        10'd63: TDATA = 39'b100000000001000100101111110110100010001;
        10'd64: TDATA = 39'b011111111111001100101111000001001100100;
        10'd65: TDATA = 39'b011111111101010100101110001011111101010;
        10'd66: TDATA = 39'b011111111011110100101101100001011011111;
        10'd67: TDATA = 39'b011111111001111100101100101100010111111;
        10'd68: TDATA = 39'b011111111000000100101011110111011010000;
        10'd69: TDATA = 39'b011111110110001100101011000010100010011;
        10'd70: TDATA = 39'b011111110100101100101010011000010100000;
        10'd71: TDATA = 39'b011111110010110100101001100011100111101;
        10'd72: TDATA = 39'b011111110000111100101000101111000001011;
        10'd73: TDATA = 39'b011111101111011100101000000101000000111;
        10'd74: TDATA = 39'b011111101101100100100111010000100101111;
        10'd75: TDATA = 39'b011111101100000100100110100110101110010;
        10'd76: TDATA = 39'b011111101010001100100101110010011110011;
        10'd77: TDATA = 39'b011111101000010100100100111110010100101;
        10'd78: TDATA = 39'b011111100110110100100100010100101010111;
        10'd79: TDATA = 39'b011111100100111100100011100000101100010;
        10'd80: TDATA = 39'b011111100011011100100010110111001011100;
        10'd81: TDATA = 39'b011111100001100100100010000011011000000;
        10'd82: TDATA = 39'b011111100000000100100001011010000000000;
        10'd83: TDATA = 39'b011111011110001100100000100110010111101;
        10'd84: TDATA = 39'b011111011100101100011111111101001000100;
        10'd85: TDATA = 39'b011111011010110100011111001001101011001;
        10'd86: TDATA = 39'b011111011001010100011110100000100100111;
        10'd87: TDATA = 39'b011111010111011100011101101101010010100;
        10'd88: TDATA = 39'b011111010101111100011101000100010101000;
        10'd89: TDATA = 39'b011111010100000100011100010001001101110;
        10'd90: TDATA = 39'b011111010010100100011011101000011001001;
        10'd91: TDATA = 39'b011111010000101100011010110101011100111;
        10'd92: TDATA = 39'b011111001111001100011010001100110001000;
        10'd93: TDATA = 39'b011111001101101100011001100100001001000;
        10'd94: TDATA = 39'b011111001011110100011000110001011100101;
        10'd95: TDATA = 39'b011111001010010100011000001000111101100;
        10'd96: TDATA = 39'b011111001000011100010111010110011100000;
        10'd97: TDATA = 39'b011111000110111100010110101110000101101;
        10'd98: TDATA = 39'b011111000101011100010110000101110011000;
        10'd99: TDATA = 39'b011111000011100100010101010011100001011;
        10'd100: TDATA = 39'b011111000010000100010100101011010111101;
        10'd101: TDATA = 39'b011111000000100100010100000011010001110;
        10'd102: TDATA = 39'b011110111110101100010011010001001111110;
        10'd103: TDATA = 39'b011110111101001100010010101001010010101;
        10'd104: TDATA = 39'b011110111011101100010010000001011001010;
        10'd105: TDATA = 39'b011110111010001100010001011001100011111;
        10'd106: TDATA = 39'b011110111000010100010000100111110110100;
        10'd107: TDATA = 39'b011110110110110100010000000000001001110;
        10'd108: TDATA = 39'b011110110101010100001111011000100000111;
        10'd109: TDATA = 39'b011110110011110100001110110000111011110;
        10'd110: TDATA = 39'b011110110001111100001101111111100010111;
        10'd111: TDATA = 39'b011110110000011100001101011000000110100;
        10'd112: TDATA = 39'b011110101110111100001100110000101110000;
        10'd113: TDATA = 39'b011110101101011100001100001001011001010;
        10'd114: TDATA = 39'b011110101011111100001011100010001000011;
        10'd115: TDATA = 39'b011110101010000100001010110001001000110;
        10'd116: TDATA = 39'b011110101000100100001010001010000000100;
        10'd117: TDATA = 39'b011110100111000100001001100010111100001;
        10'd118: TDATA = 39'b011110100101100100001000111011111011100;
        10'd119: TDATA = 39'b011110100100000100001000010100111110110;
        10'd120: TDATA = 39'b011110100010100100000111101110000101111;
        10'd121: TDATA = 39'b011110100001000100000111000111010000110;
        10'd122: TDATA = 39'b011110011111001100000110010110110011101;
        10'd123: TDATA = 39'b011110011101101100000101110000000111001;
        10'd124: TDATA = 39'b011110011100001100000101001001011110011;
        10'd125: TDATA = 39'b011110011010101100000100100010111001100;
        10'd126: TDATA = 39'b011110011001001100000011111100011000011;
        10'd127: TDATA = 39'b011110010111101100000011010101111011000;
        10'd128: TDATA = 39'b011110010110001100000010101111100001100;
        10'd129: TDATA = 39'b011110010100101100000010001001001011110;
        10'd130: TDATA = 39'b011110010011001100000001100010111001111;
        10'd131: TDATA = 39'b011110010001101100000000111100101011101;
        10'd132: TDATA = 39'b011110010000001100000000010110100001010;
        10'd133: TDATA = 39'b011110001110101011111111110000011010110;
        10'd134: TDATA = 39'b011110001101001011111111001010010111111;
        10'd135: TDATA = 39'b011110001011101011111110100100011000111;
        10'd136: TDATA = 39'b011110001010001011111101111110011101101;
        10'd137: TDATA = 39'b011110001000101011111101011000100110001;
        10'd138: TDATA = 39'b011110000111001011111100110010110010011;
        10'd139: TDATA = 39'b011110000101101011111100001101000010011;
        10'd140: TDATA = 39'b011110000100001011111011100111010110010;
        10'd141: TDATA = 39'b011110000010101011111011000001101101110;
        10'd142: TDATA = 39'b011110000001001011111010011100001001000;
        10'd143: TDATA = 39'b011101111111101011111001110110101000001;
        10'd144: TDATA = 39'b011101111110100011111001011010100001111;
        10'd145: TDATA = 39'b011101111101000011111000110101000111100;
        10'd146: TDATA = 39'b011101111011100011111000001111110000111;
        10'd147: TDATA = 39'b011101111010000011110111101010011110000;
        10'd148: TDATA = 39'b011101111000100011110111000101001110111;
        10'd149: TDATA = 39'b011101110111000011110110100000000011011;
        10'd150: TDATA = 39'b011101110101100011110101111010111011110;
        10'd151: TDATA = 39'b011101110100000011110101010101110111110;
        10'd152: TDATA = 39'b011101110010111011110100111010000111010;
        10'd153: TDATA = 39'b011101110001011011110100010101001001110;
        10'd154: TDATA = 39'b011101101111111011110011110000010000001;
        10'd155: TDATA = 39'b011101101110011011110011001011011010001;
        10'd156: TDATA = 39'b011101101100111011110010100110100111110;
        10'd157: TDATA = 39'b011101101011110011110010001011000100100;
        10'd158: TDATA = 39'b011101101010010011110001100110011000110;
        10'd159: TDATA = 39'b011101101000110011110001000001110000101;
        10'd160: TDATA = 39'b011101100111010011110000011101001100010;
        10'd161: TDATA = 39'b011101100110001011110000000001110011011;
        10'd162: TDATA = 39'b011101100100101011101111011101010101100;
        10'd163: TDATA = 39'b011101100011001011101110111000111011011;
        10'd164: TDATA = 39'b011101100001101011101110010100100100111;
        10'd165: TDATA = 39'b011101100000100011101101111001010110011;
        10'd166: TDATA = 39'b011101011111000011101101010101000110010;
        10'd167: TDATA = 39'b011101011101100011101100110000111001111;
        10'd168: TDATA = 39'b011101011100011011101100010101110011001;
        10'd169: TDATA = 39'b011101011010111011101011110001101101001;
        10'd170: TDATA = 39'b011101011001011011101011001101101010111;
        10'd171: TDATA = 39'b011101010111111011101010101001101100011;
        10'd172: TDATA = 39'b011101010110110011101010001110101111111;
        10'd173: TDATA = 39'b011101010101010011101001101010110111101;
        10'd174: TDATA = 39'b011101010100001011101001010000000000000;
        10'd175: TDATA = 39'b011101010010101011101000101100001110010;
        10'd176: TDATA = 39'b011101010001001011101000001000100000001;
        10'd177: TDATA = 39'b011101010000000011100111101101110000000;
        10'd178: TDATA = 39'b011101001110100011100111001010001000011;
        10'd179: TDATA = 39'b011101001101000011100110100110100100010;
        10'd180: TDATA = 39'b011101001011111011100110001011111011110;
        10'd181: TDATA = 39'b011101001010011011100101101000011110000;
        10'd182: TDATA = 39'b011101001001010011100101001101111010010;
        10'd183: TDATA = 39'b011101000111110011100100101010100011000;
        10'd184: TDATA = 39'b011101000110010011100100000111001111011;
        10'd185: TDATA = 39'b011101000101001011100011101100110011000;
        10'd186: TDATA = 39'b011101000011101011100011001001100101110;
        10'd187: TDATA = 39'b011101000010100011100010101111001110010;
        10'd188: TDATA = 39'b011101000001000011100010001100000111011;
        10'd189: TDATA = 39'b011100111111111011100001110001110100100;
        10'd190: TDATA = 39'b011100111110011011100001001110110100000;
        10'd191: TDATA = 39'b011100111101010011100000110100100110000;
        10'd192: TDATA = 39'b011100111011110011100000010001101011110;
        10'd193: TDATA = 39'b011100111010101011011111110111100010011;
        10'd194: TDATA = 39'b011100111001001011011111010100101110100;
        10'd195: TDATA = 39'b011100111000000011011110111010101010000;
        10'd196: TDATA = 39'b011100110110100011011110010111111100011;
        10'd197: TDATA = 39'b011100110101011011011101111101111100101;
        10'd198: TDATA = 39'b011100110011111011011101011011010101011;
        10'd199: TDATA = 39'b011100110010110011011101000001011010010;
        10'd200: TDATA = 39'b011100110001010011011100011110111001011;
        10'd201: TDATA = 39'b011100110000001011011100000101000011000;
        10'd202: TDATA = 39'b011100101111000011011011101011001110101;
        10'd203: TDATA = 39'b011100101101100011011011001000110110101;
        10'd204: TDATA = 39'b011100101100011011011010101111000111000;
        10'd205: TDATA = 39'b011100101010111011011010001100110101011;
        10'd206: TDATA = 39'b011100101001110011011001110011001010011;
        10'd207: TDATA = 39'b011100101000010011011001010000111111000;
        10'd208: TDATA = 39'b011100100111001011011000110111011000110;
        10'd209: TDATA = 39'b011100100110000011011000011101110100100;
        10'd210: TDATA = 39'b011100100100100011010111111011110010000;
        10'd211: TDATA = 39'b011100100011011011010111100010010010100;
        10'd212: TDATA = 39'b011100100010010011010111001000110101000;
        10'd213: TDATA = 39'b011100100000110011010110100110111011100;
        10'd214: TDATA = 39'b011100011111101011010110001101100010101;
        10'd215: TDATA = 39'b011100011110100011010101110100001011110;
        10'd216: TDATA = 39'b011100011101000011010101010010011011001;
        10'd217: TDATA = 39'b011100011011111011010100111001001001000;
        10'd218: TDATA = 39'b011100011010110011010100011111111000110;
        10'd219: TDATA = 39'b011100011001010011010011111110010001000;
        10'd220: TDATA = 39'b011100011000001011010011100101000101100;
        10'd221: TDATA = 39'b011100010111000011010011001011111100000;
        10'd222: TDATA = 39'b011100010101100011010010101010011101001;
        10'd223: TDATA = 39'b011100010100011011010010010001011000010;
        10'd224: TDATA = 39'b011100010011010011010001111000010101011;
        10'd225: TDATA = 39'b011100010001110011010001010110111111011;
        10'd226: TDATA = 39'b011100010000101011010000111110000001001;
        10'd227: TDATA = 39'b011100001111100011010000100101000100111;
        10'd228: TDATA = 39'b011100001110011011010000001100001010101;
        10'd229: TDATA = 39'b011100001100111011001111101011000000000;
        10'd230: TDATA = 39'b011100001011110011001111010010001010011;
        10'd231: TDATA = 39'b011100001010101011001110111001010110110;
        10'd232: TDATA = 39'b011100001001100011001110100000100101001;
        10'd233: TDATA = 39'b011100001000000011001101111111100110000;
        10'd234: TDATA = 39'b011100000110111011001101100110111001000;
        10'd235: TDATA = 39'b011100000101110011001101001110001101111;
        10'd236: TDATA = 39'b011100000100101011001100110101100100110;
        10'd237: TDATA = 39'b011100000011100011001100011100111101101;
        10'd238: TDATA = 39'b011100000010000011001011111100001100101;
        10'd239: TDATA = 39'b011100000000111011001011100011101010001;
        10'd240: TDATA = 39'b011011111111110011001011001011001001100;
        10'd241: TDATA = 39'b011011111110101011001010110010101011000;
        10'd242: TDATA = 39'b011011111101100011001010011010001110011;
        10'd243: TDATA = 39'b011011111100011011001010000001110011110;
        10'd244: TDATA = 39'b011011111010111011001001100001010011010;
        10'd245: TDATA = 39'b011011111001110011001001001000111101001;
        10'd246: TDATA = 39'b011011111000101011001000110000101001000;
        10'd247: TDATA = 39'b011011110111100011001000011000010110111;
        10'd248: TDATA = 39'b011011110110011011001000000000000110110;
        10'd249: TDATA = 39'b011011110101010011000111100111111000100;
        10'd250: TDATA = 39'b011011110100001011000111001111101100010;
        10'd251: TDATA = 39'b011011110011000011000110110111100010000;
        10'd252: TDATA = 39'b011011110001100011000110010111010111010;
        10'd253: TDATA = 39'b011011110000011011000101111111010001100;
        10'd254: TDATA = 39'b011011101111010011000101100111001101101;
        10'd255: TDATA = 39'b011011101110001011000101001111001011111;
        10'd256: TDATA = 39'b011011101101000011000100110111001011111;
        10'd257: TDATA = 39'b011011101011111011000100011111001110000;
        10'd258: TDATA = 39'b011011101010110011000100000111010010000;
        10'd259: TDATA = 39'b011011101001101011000011101111010111111;
        10'd260: TDATA = 39'b011011101000100011000011010111011111110;
        10'd261: TDATA = 39'b011011100111011011000010111111101001101;
        10'd262: TDATA = 39'b011011100110010011000010100111110101011;
        10'd263: TDATA = 39'b011011100101001011000010010000000011001;
        10'd264: TDATA = 39'b011011100100000011000001111000010010110;
        10'd265: TDATA = 39'b011011100010111011000001100000100100011;
        10'd266: TDATA = 39'b011011100001110011000001001000110111111;
        10'd267: TDATA = 39'b011011100000101011000000110001001101011;
        10'd268: TDATA = 39'b011011011111100011000000011001100100110;
        10'd269: TDATA = 39'b011011011110011011000000000001111110000;
        10'd270: TDATA = 39'b011011011101010010111111101010011001010;
        10'd271: TDATA = 39'b011011011100001010111111010010110110100;
        10'd272: TDATA = 39'b011011011011000010111110111011010101101;
        10'd273: TDATA = 39'b011011011001111010111110100011110110101;
        10'd274: TDATA = 39'b011011011000110010111110001100011001101;
        10'd275: TDATA = 39'b011011010111101010111101110100111110100;
        10'd276: TDATA = 39'b011011010110100010111101011101100101011;
        10'd277: TDATA = 39'b011011010101011010111101000110001110001;
        10'd278: TDATA = 39'b011011010100010010111100101110111000110;
        10'd279: TDATA = 39'b011011010011001010111100010111100101011;
        10'd280: TDATA = 39'b011011010010000010111100000000010011111;
        10'd281: TDATA = 39'b011011010000111010111011101001000100010;
        10'd282: TDATA = 39'b011011001111110010111011010001110110101;
        10'd283: TDATA = 39'b011011001110101010111010111010101010111;
        10'd284: TDATA = 39'b011011001101100010111010100011100001000;
        10'd285: TDATA = 39'b011011001100011010111010001100011001001;
        10'd286: TDATA = 39'b011011001011010010111001110101010011001;
        10'd287: TDATA = 39'b011011001010100010111001100101111010111;
        10'd288: TDATA = 39'b011011001001011010111001001110111000000;
        10'd289: TDATA = 39'b011011001000010010111000110111110111001;
        10'd290: TDATA = 39'b011011000111001010111000100000111000001;
        10'd291: TDATA = 39'b011011000110000010111000001001111011000;
        10'd292: TDATA = 39'b011011000100111010110111110010111111111;
        10'd293: TDATA = 39'b011011000011110010110111011100000110100;
        10'd294: TDATA = 39'b011011000010101010110111000101001111001;
        10'd295: TDATA = 39'b011011000001111010110110110110000000101;
        10'd296: TDATA = 39'b011011000000110010110110011111001100011;
        10'd297: TDATA = 39'b011010111111101010110110001000011010001;
        10'd298: TDATA = 39'b011010111110100010110101110001101001101;
        10'd299: TDATA = 39'b011010111101011010110101011010111011001;
        10'd300: TDATA = 39'b011010111100010010110101000100001110100;
        10'd301: TDATA = 39'b011010111011001010110100101101100011110;
        10'd302: TDATA = 39'b011010111010011010110100011110011101110;
        10'd303: TDATA = 39'b011010111001010010110100000111110110001;
        10'd304: TDATA = 39'b011010111000001010110011110001010000100;
        10'd305: TDATA = 39'b011010110111000010110011011010101100101;
        10'd306: TDATA = 39'b011010110101111010110011000100001010110;
        10'd307: TDATA = 39'b011010110101001010110010110101001010100;
        10'd308: TDATA = 39'b011010110100000010110010011110101011110;
        10'd309: TDATA = 39'b011010110010111010110010001000001110111;
        10'd310: TDATA = 39'b011010110001110010110001110001110011111;
        10'd311: TDATA = 39'b011010110000101010110001011011011010110;
        10'd312: TDATA = 39'b011010101111111010110001001100100000011;
        10'd313: TDATA = 39'b011010101110110010110000110110001010011;
        10'd314: TDATA = 39'b011010101101101010110000011111110110011;
        10'd315: TDATA = 39'b011010101100100010110000001001100100001;
        10'd316: TDATA = 39'b011010101011110010101111111010101110011;
        10'd317: TDATA = 39'b011010101010101010101111100100011111010;
        10'd318: TDATA = 39'b011010101001100010101111001110010010000;
        10'd319: TDATA = 39'b011010101000011010101110111000000110110;
        10'd320: TDATA = 39'b011010100111101010101110101001010101100;
        10'd321: TDATA = 39'b011010100110100010101110010011001101010;
        10'd322: TDATA = 39'b011010100101011010101101111101000110111;
        10'd323: TDATA = 39'b011010100100101010101101101110011001001;
        10'd324: TDATA = 39'b011010100011100010101101011000010101111;
        10'd325: TDATA = 39'b011010100010011010101101000010010100100;
        10'd326: TDATA = 39'b011010100001010010101100101100010101000;
        10'd327: TDATA = 39'b011010100000100010101100011101101011101;
        10'd328: TDATA = 39'b011010011111011010101100000111101111010;
        10'd329: TDATA = 39'b011010011110010010101011110001110100110;
        10'd330: TDATA = 39'b011010011101100010101011100011001110110;
        10'd331: TDATA = 39'b011010011100011010101011001101010111011;
        10'd332: TDATA = 39'b011010011011010010101010110111100001110;
        10'd333: TDATA = 39'b011010011010100010101010101000111111000;
        10'd334: TDATA = 39'b011010011001011010101010010011001100101;
        10'd335: TDATA = 39'b011010011000010010101001111101011100000;
        10'd336: TDATA = 39'b011010010111100010101001101110111100101;
        10'd337: TDATA = 39'b011010010110011010101001011001001111000;
        10'd338: TDATA = 39'b011010010101010010101001000011100011011;
        10'd339: TDATA = 39'b011010010100100010101000110101000111010;
        10'd340: TDATA = 39'b011010010011011010101000011111011110101;
        10'd341: TDATA = 39'b011010010010101010101000010001000100101;
        10'd342: TDATA = 39'b011010010001100010100111111011011111001;
        10'd343: TDATA = 39'b011010010000011010100111100101111011100;
        10'd344: TDATA = 39'b011010001111101010100111010111100100110;
        10'd345: TDATA = 39'b011010001110100010100111000010000100001;
        10'd346: TDATA = 39'b011010001101011010100110101100100101011;
        10'd347: TDATA = 39'b011010001100101010100110011110010001111;
        10'd348: TDATA = 39'b011010001011100010100110001000110110010;
        10'd349: TDATA = 39'b011010001010110010100101111010100100111;
        10'd350: TDATA = 39'b011010001001101010100101100101001100010;
        10'd351: TDATA = 39'b011010001000100010100101001111110101100;
        10'd352: TDATA = 39'b011010000111110010100101000001100111010;
        10'd353: TDATA = 39'b011010000110101010100100101100010011101;
        10'd354: TDATA = 39'b011010000101111010100100011110000111100;
        10'd355: TDATA = 39'b011010000100110010100100001000110110111;
        10'd356: TDATA = 39'b011010000100000010100011111010101100110;
        10'd357: TDATA = 39'b011010000010111010100011100101011111001;
        10'd358: TDATA = 39'b011010000001110010100011010000010011011;
        10'd359: TDATA = 39'b011010000001000010100011000010001100101;
        10'd360: TDATA = 39'b011001111111111010100010101101000011111;
        10'd361: TDATA = 39'b011001111111001010100010011110111111001;
        10'd362: TDATA = 39'b011001111110000010100010001001111001011;
        10'd363: TDATA = 39'b011001111101010010100001111011110110101;
        10'd364: TDATA = 39'b011001111100001010100001100110110100000;
        10'd365: TDATA = 39'b011001111011011010100001011000110011010;
        10'd366: TDATA = 39'b011001111010010010100001000011110011110;
        10'd367: TDATA = 39'b011001111001100010100000110101110101000;
        10'd368: TDATA = 39'b011001111000011010100000100000111000100;
        10'd369: TDATA = 39'b011001110111101010100000010010111011110;
        10'd370: TDATA = 39'b011001110110100010011111111110000010010;
        10'd371: TDATA = 39'b011001110101110010011111110000000111101;
        10'd372: TDATA = 39'b011001110100101010011111011011010001001;
        10'd373: TDATA = 39'b011001110011111010011111001101011000100;
        10'd374: TDATA = 39'b011001110010110010011110111000100101000;
        10'd375: TDATA = 39'b011001110010000010011110101010101110011;
        10'd376: TDATA = 39'b011001110000111010011110010101111101111;
        10'd377: TDATA = 39'b011001110000001010011110001000001001010;
        10'd378: TDATA = 39'b011001101111000010011101110011011011111;
        10'd379: TDATA = 39'b011001101110010010011101100101101001010;
        10'd380: TDATA = 39'b011001101101001010011101010000111110111;
        10'd381: TDATA = 39'b011001101100011010011101000011001110010;
        10'd382: TDATA = 39'b011001101011010010011100101110100110111;
        10'd383: TDATA = 39'b011001101010100010011100100000111000010;
        10'd384: TDATA = 39'b011001101001110010011100010011001010100;
        10'd385: TDATA = 39'b011001101000101010011011111110100111010;
        10'd386: TDATA = 39'b011001100111111010011011110000111011100;
        10'd387: TDATA = 39'b011001100110110010011011011100011011011;
        10'd388: TDATA = 39'b011001100110000010011011001110110001100;
        10'd389: TDATA = 39'b011001100100111010011010111010010100011;
        10'd390: TDATA = 39'b011001100100001010011010101100101100101;
        10'd391: TDATA = 39'b011001100011011010011010011111000101101;
        10'd392: TDATA = 39'b011001100010010010011010001010101100101;
        10'd393: TDATA = 39'b011001100001100010011001111101000111101;
        10'd394: TDATA = 39'b011001100000011010011001101000110001101;
        10'd395: TDATA = 39'b011001011111101010011001011011001110101;
        10'd396: TDATA = 39'b011001011110111010011001001101101100011;
        10'd397: TDATA = 39'b011001011101110010011000111001011010101;
        10'd398: TDATA = 39'b011001011101000010011000101011111010011;
        10'd399: TDATA = 39'b011001011011111010011000010111101011100;
        10'd400: TDATA = 39'b011001011011001010011000001010001101011;
        10'd401: TDATA = 39'b011001011010011010010111111100101111111;
        10'd402: TDATA = 39'b011001011001010010010111101000100101010;
        10'd403: TDATA = 39'b011001011000100010010111011011001001110;
        10'd404: TDATA = 39'b011001010111110010010111001101101111001;
        10'd405: TDATA = 39'b011001010110101010010110111001101000101;
        10'd406: TDATA = 39'b011001010101111010010110101100010000000;
        10'd407: TDATA = 39'b011001010100110010010110011000001100100;
        10'd408: TDATA = 39'b011001010100000010010110001010110101110;
        10'd409: TDATA = 39'b011001010011010010010101111101011111111;
        10'd410: TDATA = 39'b011001010010001010010101101001100000100;
        10'd411: TDATA = 39'b011001010001011010010101011100001100100;
        10'd412: TDATA = 39'b011001010000101010010101001110111001011;
        10'd413: TDATA = 39'b011001001111100010010100111010111110010;
        10'd414: TDATA = 39'b011001001110110010010100101101101101000;
        10'd415: TDATA = 39'b011001001110000010010100100000011100101;
        10'd416: TDATA = 39'b011001001100111010010100001100100101101;
        10'd417: TDATA = 39'b011001001100001010010011111111010111001;
        10'd418: TDATA = 39'b011001001011011010010011110010001001100;
        10'd419: TDATA = 39'b011001001010101010010011100100111100110;
        10'd420: TDATA = 39'b011001001001100010010011010001001011000;
        10'd421: TDATA = 39'b011001001000110010010011000100000000001;
        10'd422: TDATA = 39'b011001001000000010010010110110110110000;
        10'd423: TDATA = 39'b011001000110111010010010100011001000011;
        10'd424: TDATA = 39'b011001000110001010010010010110000000010;
        10'd425: TDATA = 39'b011001000101011010010010001000111000111;
        10'd426: TDATA = 39'b011001000100101010010001111011110010011;
        10'd427: TDATA = 39'b011001000011100010010001101000001010000;
        10'd428: TDATA = 39'b011001000010110010010001011011000101011;
        10'd429: TDATA = 39'b011001000010000010010001001110000001101;
        10'd430: TDATA = 39'b011001000000111010010000111010011101011;
        10'd431: TDATA = 39'b011001000000001010010000101101011011100;
        10'd432: TDATA = 39'b011000111111011010010000100000011010011;
        10'd433: TDATA = 39'b011000111110101010010000010011011010001;
        10'd434: TDATA = 39'b011000111101100010001111111111111011001;
        10'd435: TDATA = 39'b011000111100110010001111110010111100110;
        10'd436: TDATA = 39'b011000111100000010001111100101111111010;
        10'd437: TDATA = 39'b011000111011010010001111011001000010100;
        10'd438: TDATA = 39'b011000111010001010001111000101101000110;
        10'd439: TDATA = 39'b011000111001011010001110111000101101111;
        10'd440: TDATA = 39'b011000111000101010001110101011110011111;
        10'd441: TDATA = 39'b011000110111111010001110011110111010101;
        10'd442: TDATA = 39'b011000110111001010001110010010000010001;
        10'd443: TDATA = 39'b011000110110000010001101111110101110110;
        10'd444: TDATA = 39'b011000110101010010001101110001111000010;
        10'd445: TDATA = 39'b011000110100100010001101100101000010011;
        10'd446: TDATA = 39'b011000110011110010001101011000001101011;
        10'd447: TDATA = 39'b011000110010101010001101000100111111011;
        10'd448: TDATA = 39'b011000110001111010001100111000001100010;
        10'd449: TDATA = 39'b011000110001001010001100101011011010000;
        10'd450: TDATA = 39'b011000110000011010001100011110101000100;
        10'd451: TDATA = 39'b011000101111101010001100010001110111110;
        10'd452: TDATA = 39'b011000101110100010001011111110110000000;
        10'd453: TDATA = 39'b011000101101110010001011110010000001010;
        10'd454: TDATA = 39'b011000101101000010001011100101010011001;
        10'd455: TDATA = 39'b011000101100010010001011011000100101111;
        10'd456: TDATA = 39'b011000101011100010001011001011111001011;
        10'd457: TDATA = 39'b011000101010110010001010111111001101101;
        10'd458: TDATA = 39'b011000101001101010001010101100001101100;
        10'd459: TDATA = 39'b011000101000111010001010011111100011110;
        10'd460: TDATA = 39'b011000101000001010001010010010111010110;
        10'd461: TDATA = 39'b011000100111011010001010000110010010011;
        10'd462: TDATA = 39'b011000100110101010001001111001101010111;
        10'd463: TDATA = 39'b011000100101111010001001101101000100010;
        10'd464: TDATA = 39'b011000100100110010001001011010001011100;
        10'd465: TDATA = 39'b011000100100000010001001001101100110110;
        10'd466: TDATA = 39'b011000100011010010001001000001000010110;
        10'd467: TDATA = 39'b011000100010100010001000110100011111100;
        10'd468: TDATA = 39'b011000100001110010001000100111111100111;
        10'd469: TDATA = 39'b011000100001000010001000011011011011010;
        10'd470: TDATA = 39'b011000100000010010001000001110111010010;
        10'd471: TDATA = 39'b011000011111001010000111111100001010010;
        10'd472: TDATA = 39'b011000011110011010000111101111101011001;
        10'd473: TDATA = 39'b011000011101101010000111100011001100111;
        10'd474: TDATA = 39'b011000011100111010000111010110101111011;
        10'd475: TDATA = 39'b011000011100001010000111001010010010100;
        10'd476: TDATA = 39'b011000011011011010000110111101110110100;
        10'd477: TDATA = 39'b011000011010101010000110110001011011011;
        10'd478: TDATA = 39'b011000011001111010000110100101000000111;
        10'd479: TDATA = 39'b011000011001001010000110011000100111001;
        10'd480: TDATA = 39'b011000011000000010000110000110000010000;
        10'd481: TDATA = 39'b011000010111010010000101111001101010010;
        10'd482: TDATA = 39'b011000010110100010000101101101010011001;
        10'd483: TDATA = 39'b011000010101110010000101100000111100111;
        10'd484: TDATA = 39'b011000010101000010000101010100100111011;
        10'd485: TDATA = 39'b011000010100010010000101001000010010101;
        10'd486: TDATA = 39'b011000010011100010000100111011111110101;
        10'd487: TDATA = 39'b011000010010110010000100101111101011011;
        10'd488: TDATA = 39'b011000010010000010000100100011011000111;
        10'd489: TDATA = 39'b011000010001010010000100010111000111001;
        10'd490: TDATA = 39'b011000010000100010000100001010110110001;
        10'd491: TDATA = 39'b011000001111110010000011111110100110000;
        10'd492: TDATA = 39'b011000001111000010000011110010010110100;
        10'd493: TDATA = 39'b011000001110010010000011100110000111110;
        10'd494: TDATA = 39'b011000001101001010000011010011110011001;
        10'd495: TDATA = 39'b011000001100011010000011000111100110011;
        10'd496: TDATA = 39'b011000001011101010000010111011011010011;
        10'd497: TDATA = 39'b011000001010111010000010101111001111000;
        10'd498: TDATA = 39'b011000001010001010000010100011000100100;
        10'd499: TDATA = 39'b011000001001011010000010010110111010110;
        10'd500: TDATA = 39'b011000001000101010000010001010110001101;
        10'd501: TDATA = 39'b011000000111111010000001111110101001011;
        10'd502: TDATA = 39'b011000000111001010000001110010100001111;
        10'd503: TDATA = 39'b011000000110011010000001100110011011001;
        10'd504: TDATA = 39'b011000000101101010000001011010010101001;
        10'd505: TDATA = 39'b011000000100111010000001001110001111111;
        10'd506: TDATA = 39'b011000000100001010000001000010001011011;
        10'd507: TDATA = 39'b011000000011011010000000110110000111101;
        10'd508: TDATA = 39'b011000000010101010000000101010000100101;
        10'd509: TDATA = 39'b011000000001111010000000011110000010011;
        10'd510: TDATA = 39'b011000000001001010000000010010000000111;
        10'd511: TDATA = 39'b011000000000011010000000000110000000001;
        10'd512: TDATA = 39'b101111111110100111111111010000000001100;
        10'd513: TDATA = 39'b101111111011100111111101110000001101100;
        10'd514: TDATA = 39'b101111111000100111111100010000100101100;
        10'd515: TDATA = 39'b101111110101100111111010110001001001011;
        10'd516: TDATA = 39'b101111110010100111111001010001111001011;
        10'd517: TDATA = 39'b101111101111100111110111110010110101001;
        10'd518: TDATA = 39'b101111101100100111110110010011111101000;
        10'd519: TDATA = 39'b101111101001111111110101000001000101100;
        10'd520: TDATA = 39'b101111100110111111110011100010100011110;
        10'd521: TDATA = 39'b101111100011111111110010000100001101110;
        10'd522: TDATA = 39'b101111100000111111110000100110000011101;
        10'd523: TDATA = 39'b101111011110010111101111010011110100101;
        10'd524: TDATA = 39'b101111011011010111101101110110000000110;
        10'd525: TDATA = 39'b101111011000010111101100011000011000111;
        10'd526: TDATA = 39'b101111010101010111101010111010111100110;
        10'd527: TDATA = 39'b101111010010101111101001101001010101111;
        10'd528: TDATA = 39'b101111001111101111101000001100001111111;
        10'd529: TDATA = 39'b101111001100101111100110101111010101110;
        10'd530: TDATA = 39'b101111001010000111100101011110001100101;
        10'd531: TDATA = 39'b101111000111000111100100000001101000101;
        10'd532: TDATA = 39'b101111000100011111100010110000110010110;
        10'd533: TDATA = 39'b101111000001011111100001010100100100111;
        10'd534: TDATA = 39'b101110111110110111100000000100000010010;
        10'd535: TDATA = 39'b101110111011110111011110101000001010011;
        10'd536: TDATA = 39'b101110111001001111011101010111111011001;
        10'd537: TDATA = 39'b101110110110001111011011111100011001001;
        10'd538: TDATA = 39'b101110110011100111011010101100011101001;
        10'd539: TDATA = 39'b101110110000100111011001010001010001001;
        10'd540: TDATA = 39'b101110101101111111011000000001101000010;
        10'd541: TDATA = 39'b101110101011010111010110110010001000011;
        10'd542: TDATA = 39'b101110101000010111010101010111011100100;
        10'd543: TDATA = 39'b101110100101101111010100001000001111110;
        10'd544: TDATA = 39'b101110100011000111010010111001001011111;
        10'd545: TDATA = 39'b101110100000000111010001011111000000000;
        10'd546: TDATA = 39'b101110011101011111010000010000001111010;
        10'd547: TDATA = 39'b101110011010110111001111000001100111010;
        10'd548: TDATA = 39'b101110011000001111001101110011001000010;
        10'd549: TDATA = 39'b101110010101100111001100100100110010001;
        10'd550: TDATA = 39'b101110010010100111001011001011011010100;
        10'd551: TDATA = 39'b101110001111111111001001111101010111011;
        10'd552: TDATA = 39'b101110001101010111001000101111011101001;
        10'd553: TDATA = 39'b101110001010101111000111100001101011101;
        10'd554: TDATA = 39'b101110001000000111000110010100000011000;
        10'd555: TDATA = 39'b101110000101011111000101000110100011010;
        10'd556: TDATA = 39'b101110000010110111000011111001001100010;
        10'd557: TDATA = 39'b101110000000001111000010101011111110001;
        10'd558: TDATA = 39'b101101111101100111000001011110111000110;
        10'd559: TDATA = 39'b101101111010111111000000010001111100001;
        10'd560: TDATA = 39'b101101111000010110111111000101001000011;
        10'd561: TDATA = 39'b101101110101101110111101111000011101011;
        10'd562: TDATA = 39'b101101110011000110111100101011111011010;
        10'd563: TDATA = 39'b101101110000011110111011011111100001110;
        10'd564: TDATA = 39'b101101101101110110111010010011010001001;
        10'd565: TDATA = 39'b101101101011001110111001000111001001001;
        10'd566: TDATA = 39'b101101101000100110110111111011001010000;
        10'd567: TDATA = 39'b101101100101111110110110101111010011100;
        10'd568: TDATA = 39'b101101100011010110110101100011100101110;
        10'd569: TDATA = 39'b101101100000101110110100011000000000110;
        10'd570: TDATA = 39'b101101011110011110110011010111010101101;
        10'd571: TDATA = 39'b101101011011110110110010001100000000111;
        10'd572: TDATA = 39'b101101011001001110110001000000110100110;
        10'd573: TDATA = 39'b101101010110100110101111110101110001010;
        10'd574: TDATA = 39'b101101010100010110101110110101100010111;
        10'd575: TDATA = 39'b101101010001101110101101101010101111100;
        10'd576: TDATA = 39'b101101001111000110101100100000000100111;
        10'd577: TDATA = 39'b101101001100011110101011010101100010111;
        10'd578: TDATA = 39'b101101001010001110101010010101110001001;
        10'd579: TDATA = 39'b101101000111100110101001001011011111001;
        10'd580: TDATA = 39'b101101000100111110101000000001010101111;
        10'd581: TDATA = 39'b101101000010101110100111000001111001010;
        10'd582: TDATA = 39'b101101000000000110100101111000000000000;
        10'd583: TDATA = 39'b101100111101110110100100111000110001001;
        10'd584: TDATA = 39'b101100111011001110100011101111000111111;
        10'd585: TDATA = 39'b101100111000111110100010110000000110110;
        10'd586: TDATA = 39'b101100110110010110100001100110101101011;
        10'd587: TDATA = 39'b101100110100000110100000100111111001111;
        10'd588: TDATA = 39'b101100110001011110011111011110110000100;
        10'd589: TDATA = 39'b101100101111001110011110100000001010101;
        10'd590: TDATA = 39'b101100101100100110011101010111010001001;
        10'd591: TDATA = 39'b101100101010010110011100011000111000111;
        10'd592: TDATA = 39'b101100100111101110011011010000001111010;
        10'd593: TDATA = 39'b101100100101011110011010010010000100110;
        10'd594: TDATA = 39'b101100100010110110011001001001101010111;
        10'd595: TDATA = 39'b101100100000100110011000001011101101111;
        10'd596: TDATA = 39'b101100011110010110010111001101110111001;
        10'd597: TDATA = 39'b101100011011101110010110000101110100100;
        10'd598: TDATA = 39'b101100011001011110010101001000001011010;
        10'd599: TDATA = 39'b101100010111001110010100001010101000010;
        10'd600: TDATA = 39'b101100010100100110010011000010111100110;
        10'd601: TDATA = 39'b101100010010010110010010000101100111010;
        10'd602: TDATA = 39'b101100010000000110010001001000011000000;
        10'd603: TDATA = 39'b101100001101011110010000000001000011011;
        10'd604: TDATA = 39'b101100001011001110001111000100000001101;
        10'd605: TDATA = 39'b101100001000111110001110000111000110001;
        10'd606: TDATA = 39'b101100000110101110001101001010010000110;
        10'd607: TDATA = 39'b101100000100011110001100001101100001101;
        10'd608: TDATA = 39'b101100000001110110001011000110110010100;
        10'd609: TDATA = 39'b101011111111100110001010001010010000110;
        10'd610: TDATA = 39'b101011111101010110001001001101110101010;
        10'd611: TDATA = 39'b101011111011000110001000010001011111111;
        10'd612: TDATA = 39'b101011111000110110000111010101010000101;
        10'd613: TDATA = 39'b101011110110100110000110011001000111101;
        10'd614: TDATA = 39'b101011110100010110000101011101000100111;
        10'd615: TDATA = 39'b101011110010000110000100100001001000001;
        10'd616: TDATA = 39'b101011101111011110000011011011010011111;
        10'd617: TDATA = 39'b101011101101001110000010011111100100100;
        10'd618: TDATA = 39'b101011101010111110000001100011111011010;
        10'd619: TDATA = 39'b101011101000101110000000101000011000010;
        10'd620: TDATA = 39'b101011100110011101111111101100111011011;
        10'd621: TDATA = 39'b101011100100001101111110110001100100100;
        10'd622: TDATA = 39'b101011100001111101111101110110010011111;
        10'd623: TDATA = 39'b101011011111101101111100111011001001011;
        10'd624: TDATA = 39'b101011011101110101111100001001111010100;
        10'd625: TDATA = 39'b101011011011100101111011001110111011010;
        10'd626: TDATA = 39'b101011011001010101111010010100000010000;
        10'd627: TDATA = 39'b101011010111000101111001011001001110111;
        10'd628: TDATA = 39'b101011010100110101111000011110100001111;
        10'd629: TDATA = 39'b101011010010100101110111100011111010111;
        10'd630: TDATA = 39'b101011010000010101110110101001011010001;
        10'd631: TDATA = 39'b101011001110000101110101101110111111011;
        10'd632: TDATA = 39'b101011001011110101110100110100101010101;
        10'd633: TDATA = 39'b101011001001111101110100000100001000110;
        10'd634: TDATA = 39'b101011000111101101110011001001111111001;
        10'd635: TDATA = 39'b101011000101011101110010001111111011101;
        10'd636: TDATA = 39'b101011000011001101110001010101111110010;
        10'd637: TDATA = 39'b101011000001010101110000100101101111101;
        10'd638: TDATA = 39'b101010111111000101101111101011111101011;
        10'd639: TDATA = 39'b101010111100110101101110110010010001000;
        10'd640: TDATA = 39'b101010111010100101101101111000101010110;
        10'd641: TDATA = 39'b101010111000101101101101001000101111100;
        10'd642: TDATA = 39'b101010110110011101101100001111010100011;
        10'd643: TDATA = 39'b101010110100001101101011010101111111001;
        10'd644: TDATA = 39'b101010110010010101101010100110010010001;
        10'd645: TDATA = 39'b101010110000000101101001101101001000000;
        10'd646: TDATA = 39'b101010101101110101101000110100000011111;
        10'd647: TDATA = 39'b101010101011111101101000000100100101000;
        10'd648: TDATA = 39'b101010101001101101100111001011101011111;
        10'd649: TDATA = 39'b101010100111011101100110010010111000110;
        10'd650: TDATA = 39'b101010100101100101100101100011101000001;
        10'd651: TDATA = 39'b101010100011010101100100101011000000000;
        10'd652: TDATA = 39'b101010100001011101100011111011111000100;
        10'd653: TDATA = 39'b101010011111001101100011000011011011010;
        10'd654: TDATA = 39'b101010011101010101100010010100011100111;
        10'd655: TDATA = 39'b101010011011000101100001011100001010101;
        10'd656: TDATA = 39'b101010011000110101100000100011111110011;
        10'd657: TDATA = 39'b101010010110111101011111110101001110001;
        10'd658: TDATA = 39'b101010010100101101011110111101001100110;
        10'd659: TDATA = 39'b101010010010110101011110001110100101100;
        10'd660: TDATA = 39'b101010010000111101011101100000000010100;
        10'd661: TDATA = 39'b101010001110101101011100101000010001000;
        10'd662: TDATA = 39'b101010001100110101011011111001110111000;
        10'd663: TDATA = 39'b101010001010100101011011000010010000011;
        10'd664: TDATA = 39'b101010001000101101011010010011111111100;
        10'd665: TDATA = 39'b101010000110011101011001011100100011110;
        10'd666: TDATA = 39'b101010000100100101011000101110011011111;
        10'd667: TDATA = 39'b101010000010101101011000000000011000000;
        10'd668: TDATA = 39'b101010000000011101010111001001001100001;
        10'd669: TDATA = 39'b101001111110100101010110011011010001010;
        10'd670: TDATA = 39'b101001111100101101010101101101011010101;
        10'd671: TDATA = 39'b101001111010011101010100110110011110100;
        10'd672: TDATA = 39'b101001111000100101010100001000110000110;
        10'd673: TDATA = 39'b101001110110101101010011011011000111010;
        10'd674: TDATA = 39'b101001110100011101010010100100011010110;
        10'd675: TDATA = 39'b101001110010100101010001110110111010001;
        10'd676: TDATA = 39'b101001110000101101010001001001011101101;
        10'd677: TDATA = 39'b101001101110011101010000010011000000110;
        10'd678: TDATA = 39'b101001101100100101001111100101101101010;
        10'd679: TDATA = 39'b101001101010101101001110111000011101111;
        10'd680: TDATA = 39'b101001101000110101001110001011010010011;
        10'd681: TDATA = 39'b101001100110111101001101011110001011001;
        10'd682: TDATA = 39'b101001100100101101001100101000000111101;
        10'd683: TDATA = 39'b101001100010110101001011111011001001010;
        10'd684: TDATA = 39'b101001100000111101001011001110001110111;
        10'd685: TDATA = 39'b101001011111000101001010100001011000101;
        10'd686: TDATA = 39'b101001011101001101001001110100100110011;
        10'd687: TDATA = 39'b101001011010111101001000111110111100010;
        10'd688: TDATA = 39'b101001011001000101001000010010010011000;
        10'd689: TDATA = 39'b101001010111001101000111100101101101101;
        10'd690: TDATA = 39'b101001010101010101000110111001001100011;
        10'd691: TDATA = 39'b101001010011011101000110001100101111010;
        10'd692: TDATA = 39'b101001010001100101000101100000010110000;
        10'd693: TDATA = 39'b101001001111101101000100110100000000111;
        10'd694: TDATA = 39'b101001001101110101000100000111101111110;
        10'd695: TDATA = 39'b101001001011111101000011011011100010101;
        10'd696: TDATA = 39'b101001001010000101000010101111011001101;
        10'd697: TDATA = 39'b101001001000001101000010000011010100100;
        10'd698: TDATA = 39'b101001000110010101000001010111010011100;
        10'd699: TDATA = 39'b101001000100011101000000101011010110100;
        10'd700: TDATA = 39'b101001000010100100111111111111011101100;
        10'd701: TDATA = 39'b101001000000101100111111010011101000100;
        10'd702: TDATA = 39'b101000111110110100111110100111110111100;
        10'd703: TDATA = 39'b101000111100111100111101111100001010100;
        10'd704: TDATA = 39'b101000111011000100111101010000100001100;
        10'd705: TDATA = 39'b101000111001001100111100100100111100100;
        10'd706: TDATA = 39'b101000110111010100111011111001011011100;
        10'd707: TDATA = 39'b101000110101011100111011001101111110100;
        10'd708: TDATA = 39'b101000110011100100111010100010100101011;
        10'd709: TDATA = 39'b101000110001101100111001110111010000011;
        10'd710: TDATA = 39'b101000101111110100111001001011111111011;
        10'd711: TDATA = 39'b101000101101111100111000100000110010010;
        10'd712: TDATA = 39'b101000101100000100110111110101101001001;
        10'd713: TDATA = 39'b101000101010001100110111001010100100000;
        10'd714: TDATA = 39'b101000101000101100110110101000001001001;
        10'd715: TDATA = 39'b101000100110110100110101111101001011001;
        10'd716: TDATA = 39'b101000100100111100110101010010010001001;
        10'd717: TDATA = 39'b101000100011000100110100100111011011001;
        10'd718: TDATA = 39'b101000100001001100110011111100101001000;
        10'd719: TDATA = 39'b101000011111101100110011011010011101011;
        10'd720: TDATA = 39'b101000011101110100110010101111110010011;
        10'd721: TDATA = 39'b101000011011111100110010000101001011011;
        10'd722: TDATA = 39'b101000011010000100110001011010101000010;
        10'd723: TDATA = 39'b101000011000001100110000110000001001001;
        10'd724: TDATA = 39'b101000010110101100110000001110001100101;
        10'd725: TDATA = 39'b101000010100110100101111100011110100101;
        10'd726: TDATA = 39'b101000010010111100101110111001100000100;
        10'd727: TDATA = 39'b101000010001000100101110001111010000011;
        10'd728: TDATA = 39'b101000001111100100101101101101011111111;
        10'd729: TDATA = 39'b101000001101101100101101000011010110110;
        10'd730: TDATA = 39'b101000001011110100101100011001010001100;
        10'd731: TDATA = 39'b101000001010010100101011110111101001111;
        10'd732: TDATA = 39'b101000001000011100101011001101101011110;
        10'd733: TDATA = 39'b101000000110100100101010100011110001101;
        10'd734: TDATA = 39'b101000000101000100101010000010010010101;
        10'd735: TDATA = 39'b101000000011001100101001011000011111100;
        10'd736: TDATA = 39'b101000000001010100101000101110110000010;
        10'd737: TDATA = 39'b100111111111110100101000001101011010001;
        10'd738: TDATA = 39'b100111111101111100100111100011110001111;
        10'd739: TDATA = 39'b100111111100000100100110111010001101101;
        10'd740: TDATA = 39'b100111111010100100100110011001000000010;
        10'd741: TDATA = 39'b100111111000101100100101101111100010111;
        10'd742: TDATA = 39'b100111110111001100100101001110011011001;
        10'd743: TDATA = 39'b100111110101010100100100100101000100111;
        10'd744: TDATA = 39'b100111110011011100100011111011110010100;
        10'd745: TDATA = 39'b100111110001111100100011011010110011011;
        10'd746: TDATA = 39'b100111110000000100100010110001101000000;
        10'd747: TDATA = 39'b100111101110100100100010010000101110100;
        10'd748: TDATA = 39'b100111101100101100100001100111101010001;
        10'd749: TDATA = 39'b100111101011001100100001000110110110001;
        10'd750: TDATA = 39'b100111101001010100100000011101111000110;
        10'd751: TDATA = 39'b100111100111110100011111111101001010011;
        10'd752: TDATA = 39'b100111100101111100011111010100010100000;
        10'd753: TDATA = 39'b100111100100011100011110110011101011001;
        10'd754: TDATA = 39'b100111100010100100011110001010111011110;
        10'd755: TDATA = 39'b100111100001000100011101101010011000100;
        10'd756: TDATA = 39'b100111011111001100011101000001101111111;
        10'd757: TDATA = 39'b100111011101101100011100100001010010010;
        10'd758: TDATA = 39'b100111011011110100011011111000110000101;
        10'd759: TDATA = 39'b100111011010010100011011011000011000100;
        10'd760: TDATA = 39'b100111011000110100011010111000000010111;
        10'd761: TDATA = 39'b100111010110111100011010001111101011010;
        10'd762: TDATA = 39'b100111010101011100011001101111011011010;
        10'd763: TDATA = 39'b100111010011100100011001000111001010100;
        10'd764: TDATA = 39'b100111010010000100011000100110111111111;
        10'd765: TDATA = 39'b100111010000100100011000000110110111110;
        10'd766: TDATA = 39'b100111001110101100010111011110110001001;
        10'd767: TDATA = 39'b100111001101001100010110111110101110100;
        10'd768: TDATA = 39'b100111001011101100010110011110101110011;
        10'd769: TDATA = 39'b100111001001110100010101110110110001100;
        10'd770: TDATA = 39'b100111001000010100010101010110110110111;
        10'd771: TDATA = 39'b100111000110110100010100110110111110110;
        10'd772: TDATA = 39'b100111000100111100010100001111001011111;
        10'd773: TDATA = 39'b100111000011011100010011101111011001001;
        10'd774: TDATA = 39'b100111000001111100010011001111101000111;
        10'd775: TDATA = 39'b100111000000000100010010101000000000000;
        10'd776: TDATA = 39'b100110111110100100010010001000010101010;
        10'd777: TDATA = 39'b100110111101000100010001101000101100111;
        10'd778: TDATA = 39'b100110111011001100010001000001001101111;
        10'd779: TDATA = 39'b100110111001101100010000100001101011000;
        10'd780: TDATA = 39'b100110111000001100010000000010001010100;
        10'd781: TDATA = 39'b100110110110101100001111100010101100100;
        10'd782: TDATA = 39'b100110110100110100001110111011011010100;
        10'd783: TDATA = 39'b100110110011010100001110011100000001111;
        10'd784: TDATA = 39'b100110110001110100001101111100101011110;
        10'd785: TDATA = 39'b100110110000010100001101011101011000001;
        10'd786: TDATA = 39'b100110101110110100001100111110000110110;
        10'd787: TDATA = 39'b100110101100111100001100010111000100101;
        10'd788: TDATA = 39'b100110101011011100001011110111111000110;
        10'd789: TDATA = 39'b100110101001111100001011011000101111011;
        10'd790: TDATA = 39'b100110101000011100001010111001101000011;
        10'd791: TDATA = 39'b100110100110111100001010011010100011110;
        10'd792: TDATA = 39'b100110100101011100001001111011100001101;
        10'd793: TDATA = 39'b100110100011100100001001010100110010010;
        10'd794: TDATA = 39'b100110100010000100001000110101110101100;
        10'd795: TDATA = 39'b100110100000100100001000010110111011010;
        10'd796: TDATA = 39'b100110011111000100000111111000000011010;
        10'd797: TDATA = 39'b100110011101100100000111011001001101110;
        10'd798: TDATA = 39'b100110011100000100000110111010011010101;
        10'd799: TDATA = 39'b100110011010100100000110011011101001111;
        10'd800: TDATA = 39'b100110011001000100000101111100111011101;
        10'd801: TDATA = 39'b100110010111001100000101010110100101000;
        10'd802: TDATA = 39'b100110010101101100000100110111111100001;
        10'd803: TDATA = 39'b100110010100001100000100011001010101101;
        10'd804: TDATA = 39'b100110010010101100000011111010110001100;
        10'd805: TDATA = 39'b100110010001001100000011011100001111110;
        10'd806: TDATA = 39'b100110001111101100000010111101110000011;
        10'd807: TDATA = 39'b100110001110001100000010011111010011011;
        10'd808: TDATA = 39'b100110001100101100000010000000111000111;
        10'd809: TDATA = 39'b100110001011001100000001100010100000101;
        10'd810: TDATA = 39'b100110001001101100000001000100001010111;
        10'd811: TDATA = 39'b100110001000001100000000100101110111100;
        10'd812: TDATA = 39'b100110000110101100000000000111100110100;
        10'd813: TDATA = 39'b100110000101001011111111101001010111110;
        10'd814: TDATA = 39'b100110000011101011111111001011001011100;
        10'd815: TDATA = 39'b100110000010001011111110101101000001101;
        10'd816: TDATA = 39'b100110000000101011111110001110111010001;
        10'd817: TDATA = 39'b100101111111001011111101110000110101000;
        10'd818: TDATA = 39'b100101111101101011111101010010110010010;
        10'd819: TDATA = 39'b100101111100001011111100110100110001111;
        10'd820: TDATA = 39'b100101111010101011111100010110110011111;
        10'd821: TDATA = 39'b100101111001001011111011111000111000001;
        10'd822: TDATA = 39'b100101110111101011111011011010111110111;
        10'd823: TDATA = 39'b100101110110001011111010111101001000000;
        10'd824: TDATA = 39'b100101110100101011111010011111010011100;
        10'd825: TDATA = 39'b100101110011100011111010001000111101101;
        10'd826: TDATA = 39'b100101110010000011111001101011001101001;
        10'd827: TDATA = 39'b100101110000100011111001001101011111001;
        10'd828: TDATA = 39'b100101101111000011111000101111110011011;
        10'd829: TDATA = 39'b100101101101100011111000010010001010001;
        10'd830: TDATA = 39'b100101101100000011110111110100100011001;
        10'd831: TDATA = 39'b100101101010100011110111010110111110100;
        10'd832: TDATA = 39'b100101101001000011110110111001011100010;
        10'd833: TDATA = 39'b100101100111111011110110100011010100001;
        10'd834: TDATA = 39'b100101100110011011110110000101110101111;
        10'd835: TDATA = 39'b100101100100111011110101101000011010001;
        10'd836: TDATA = 39'b100101100011011011110101001011000000101;
        10'd837: TDATA = 39'b100101100001111011110100101101101001101;
        10'd838: TDATA = 39'b100101100000011011110100010000010100111;
        10'd839: TDATA = 39'b100101011111010011110011111010010110110;
        10'd840: TDATA = 39'b100101011101110011110011011101000110001;
        10'd841: TDATA = 39'b100101011100010011110010111111110111111;
        10'd842: TDATA = 39'b100101011010110011110010100010101011111;
        10'd843: TDATA = 39'b100101011001010011110010000101100010010;
        10'd844: TDATA = 39'b100101011000001011110001101111101100100;
        10'd845: TDATA = 39'b100101010110101011110001010010100111000;
        10'd846: TDATA = 39'b100101010101001011110000110101100011110;
        10'd847: TDATA = 39'b100101010011101011110000011000100010111;
        10'd848: TDATA = 39'b100101010010100011110000000010110011110;
        10'd849: TDATA = 39'b100101010001000011101111100101110111000;
        10'd850: TDATA = 39'b100101001111100011101111001000111100100;
        10'd851: TDATA = 39'b100101001110000011101110101100000100011;
        10'd852: TDATA = 39'b100101001100111011101110010110011011110;
        10'd853: TDATA = 39'b100101001011011011101101111001100111101;
        10'd854: TDATA = 39'b100101001001111011101101011100110101111;
        10'd855: TDATA = 39'b100101001000011011101101000000000110100;
        10'd856: TDATA = 39'b100101000111010011101100101010100100100;
        10'd857: TDATA = 39'b100101000101110011101100001101111001001;
        10'd858: TDATA = 39'b100101000100010011101011110001010000000;
        10'd859: TDATA = 39'b100101000011001011101011011011110010110;
        10'd860: TDATA = 39'b100101000001101011101010111111001101110;
        10'd861: TDATA = 39'b100101000000001011101010100010101011001;
        10'd862: TDATA = 39'b100100111111000011101010001101010010101;
        10'd863: TDATA = 39'b100100111101100011101001110000110100000;
        10'd864: TDATA = 39'b100100111100000011101001010100010111101;
        10'd865: TDATA = 39'b100100111010111011101000111111000011111;
        10'd866: TDATA = 39'b100100111001011011101000100010101011101;
        10'd867: TDATA = 39'b100100110111111011101000000110010101101;
        10'd868: TDATA = 39'b100100110110110011100111110001000110101;
        10'd869: TDATA = 39'b100100110101010011100111010100110100110;
        10'd870: TDATA = 39'b100100110100001011100110111111101000110;
        10'd871: TDATA = 39'b100100110010101011100110100011011010111;
        10'd872: TDATA = 39'b100100110001001011100110000111001111010;
        10'd873: TDATA = 39'b100100110000000011100101110010001000000;
        10'd874: TDATA = 39'b100100101110100011100101010110000000011;
        10'd875: TDATA = 39'b100100101101011011100101000000111100010;
        10'd876: TDATA = 39'b100100101011111011100100100100111000101;
        10'd877: TDATA = 39'b100100101010110011100100001111110111011;
        10'd878: TDATA = 39'b100100101001010011100011110011110111111;
        10'd879: TDATA = 39'b100100100111110011100011010111111010101;
        10'd880: TDATA = 39'b100100100110101011100011000010111110001;
        10'd881: TDATA = 39'b100100100101001011100010100111000100111;
        10'd882: TDATA = 39'b100100100100000011100010010010001011011;
        10'd883: TDATA = 39'b100100100010100011100001110110010110001;
        10'd884: TDATA = 39'b100100100001011011100001100001011111101;
        10'd885: TDATA = 39'b100100011111111011100001000101101110011;
        10'd886: TDATA = 39'b100100011110110011100000110000111010111;
        10'd887: TDATA = 39'b100100011101010011100000010101001101101;
        10'd888: TDATA = 39'b100100011100001011100000000000011101001;
        10'd889: TDATA = 39'b100100011010101011011111100100110011110;
        10'd890: TDATA = 39'b100100011001100011011111010000000110011;
        10'd891: TDATA = 39'b100100011000000011011110110100100001000;
        10'd892: TDATA = 39'b100100010110111011011110011111110110100;
        10'd893: TDATA = 39'b100100010101011011011110000100010101001;
        10'd894: TDATA = 39'b100100010100010011011101101111101101101;
        10'd895: TDATA = 39'b100100010010110011011101010100010000010;
        10'd896: TDATA = 39'b100100010001101011011100111111101011110;
        10'd897: TDATA = 39'b100100010000001011011100100100010010010;
        10'd898: TDATA = 39'b100100001111000011011100001111110000110;
        10'd899: TDATA = 39'b100100001101111011011011111011010000100;
        10'd900: TDATA = 39'b100100001100011011011011011111111100110;
        10'd901: TDATA = 39'b100100001011010011011011001011011111011;
        10'd902: TDATA = 39'b100100001001110011011010110000001111101;
        10'd903: TDATA = 39'b100100001000101011011010011011110101010;
        10'd904: TDATA = 39'b100100000111001011011010000000101001011;
        10'd905: TDATA = 39'b100100000110000011011001101100010010000;
        10'd906: TDATA = 39'b100100000100111011011001010111111011111;
        10'd907: TDATA = 39'b100100000011011011011000111100110101110;
        10'd908: TDATA = 39'b100100000010010011011000101000100010100;
        10'd909: TDATA = 39'b100100000000110011011000001101100000010;
        10'd910: TDATA = 39'b100011111111101011010111111001010000001;
        10'd911: TDATA = 39'b100011111110100011010111100101000001001;
        10'd912: TDATA = 39'b100011111101000011010111001010000100100;
        10'd913: TDATA = 39'b100011111011111011010110110101111000100;
        10'd914: TDATA = 39'b100011111010110011010110100001101101110;
        10'd915: TDATA = 39'b100011111001010011010110000110110110110;
        10'd916: TDATA = 39'b100011111000001011010101110010101111000;
        10'd917: TDATA = 39'b100011110111000011010101011110101000100;
        10'd918: TDATA = 39'b100011110101100011010101000011110111000;
        10'd919: TDATA = 39'b100011110100011011010100101111110011100;
        10'd920: TDATA = 39'b100011110011010011010100011011110001001;
        10'd921: TDATA = 39'b100011110001110011010100000001000101011;
        10'd922: TDATA = 39'b100011110000101011010011101101000101111;
        10'd923: TDATA = 39'b100011101111100011010011011001000111110;
        10'd924: TDATA = 39'b100011101110000011010010111110100001101;
        10'd925: TDATA = 39'b100011101100111011010010101010100110011;
        10'd926: TDATA = 39'b100011101011110011010010010110101100011;
        10'd927: TDATA = 39'b100011101010101011010010000010110011110;
        10'd928: TDATA = 39'b100011101001001011010001101000010100110;
        10'd929: TDATA = 39'b100011101000000011010001010100011111000;
        10'd930: TDATA = 39'b100011100110111011010001000000101010100;
        10'd931: TDATA = 39'b100011100101011011010000100110010001001;
        10'd932: TDATA = 39'b100011100100010011010000010010011111100;
        10'd933: TDATA = 39'b100011100011001011001111111110101111001;
        10'd934: TDATA = 39'b100011100010000011001111101011000000000;
        10'd935: TDATA = 39'b100011100000100011001111010000101101111;
        10'd936: TDATA = 39'b100011011111011011001110111101000001101;
        10'd937: TDATA = 39'b100011011110010011001110101001010110110;
        10'd938: TDATA = 39'b100011011101001011001110010101101101001;
        10'd939: TDATA = 39'b100011011100000011001110000010000100101;
        10'd940: TDATA = 39'b100011011010100011001101100111111011010;
        10'd941: TDATA = 39'b100011011001011011001101010100010101110;
        10'd942: TDATA = 39'b100011011000010011001101000000110001100;
        10'd943: TDATA = 39'b100011010111001011001100101101001110100;
        10'd944: TDATA = 39'b100011010101101011001100010011001100011;
        10'd945: TDATA = 39'b100011010100100011001011111111101100001;
        10'd946: TDATA = 39'b100011010011011011001011101100001101010;
        10'd947: TDATA = 39'b100011010010010011001011011000101111101;
        10'd948: TDATA = 39'b100011010001001011001011000101010011001;
        10'd949: TDATA = 39'b100011010000000011001010110001111000000;
        10'd950: TDATA = 39'b100011001110100011001010011000000000011;
        10'd951: TDATA = 39'b100011001101011011001010000100101000000;
        10'd952: TDATA = 39'b100011001100010011001001110001010001000;
        10'd953: TDATA = 39'b100011001011001011001001011101111011010;
        10'd954: TDATA = 39'b100011001010000011001001001010100110101;
        10'd955: TDATA = 39'b100011001000111011001000110111010011010;
        10'd956: TDATA = 39'b100011000111110011001000100100000001001;
        10'd957: TDATA = 39'b100011000110010011001000001010010101101;
        10'd958: TDATA = 39'b100011000101001011000111110111000110011;
        10'd959: TDATA = 39'b100011000100000011000111100011111000011;
        10'd960: TDATA = 39'b100011000010111011000111010000101011101;
        10'd961: TDATA = 39'b100011000001110011000110111101100000001;
        10'd962: TDATA = 39'b100011000000101011000110101010010101110;
        10'd963: TDATA = 39'b100010111111100011000110010111001100110;
        10'd964: TDATA = 39'b100010111110011011000110000100000100111;
        10'd965: TDATA = 39'b100010111101010011000101110000111110010;
        10'd966: TDATA = 39'b100010111011110011000101010111100010000;
        10'd967: TDATA = 39'b100010111010101011000101000100011110010;
        10'd968: TDATA = 39'b100010111001100011000100110001011011110;
        10'd969: TDATA = 39'b100010111000011011000100011110011010100;
        10'd970: TDATA = 39'b100010110111010011000100001011011010011;
        10'd971: TDATA = 39'b100010110110001011000011111000011011101;
        10'd972: TDATA = 39'b100010110101000011000011100101011110000;
        10'd973: TDATA = 39'b100010110011111011000011010010100001101;
        10'd974: TDATA = 39'b100010110010110011000010111111100110011;
        10'd975: TDATA = 39'b100010110001101011000010101100101100100;
        10'd976: TDATA = 39'b100010110000100011000010011001110011110;
        10'd977: TDATA = 39'b100010101111011011000010000110111100010;
        10'd978: TDATA = 39'b100010101110010011000001110100000110000;
        10'd979: TDATA = 39'b100010101101001011000001100001010001000;
        10'd980: TDATA = 39'b100010101100000011000001001110011101001;
        10'd981: TDATA = 39'b100010101010111011000000111011101010100;
        10'd982: TDATA = 39'b100010101001110011000000101000111001001;
        10'd983: TDATA = 39'b100010101000101011000000010110001001000;
        10'd984: TDATA = 39'b100010100111100011000000000011011010000;
        10'd985: TDATA = 39'b100010100110011010111111110000101100010;
        10'd986: TDATA = 39'b100010100101010010111111011101111111110;
        10'd987: TDATA = 39'b100010100100001010111111001011010100011;
        10'd988: TDATA = 39'b100010100011000010111110111000101010011;
        10'd989: TDATA = 39'b100010100001111010111110100110000001011;
        10'd990: TDATA = 39'b100010100000110010111110010011011001110;
        10'd991: TDATA = 39'b100010011111101010111110000000110011011;
        10'd992: TDATA = 39'b100010011110100010111101101110001110001;
        10'd993: TDATA = 39'b100010011101011010111101011011101010000;
        10'd994: TDATA = 39'b100010011100010010111101001001000111010;
        10'd995: TDATA = 39'b100010011011001010111100110110100101101;
        10'd996: TDATA = 39'b100010011010000010111100100100000101010;
        10'd997: TDATA = 39'b100010011000111010111100010001100110000;
        10'd998: TDATA = 39'b100010010111110010111011111111001000001;
        10'd999: TDATA = 39'b100010010110101010111011101100101011010;
        10'd1000: TDATA = 39'b100010010101100010111011011010001111110;
        10'd1001: TDATA = 39'b100010010100011010111011000111110101011;
        10'd1002: TDATA = 39'b100010010011010010111010110101011100010;
        10'd1003: TDATA = 39'b100010010010001010111010100011000100010;
        10'd1004: TDATA = 39'b100010010001011010111010010110110101000;
        10'd1005: TDATA = 39'b100010010000010010111010000100011111001;
        10'd1006: TDATA = 39'b100010001111001010111001110010001010011;
        10'd1007: TDATA = 39'b100010001110000010111001011111110110111;
        10'd1008: TDATA = 39'b100010001100111010111001001101100100100;
        10'd1009: TDATA = 39'b100010001011110010111000111011010011011;
        10'd1010: TDATA = 39'b100010001010101010111000101001000011100;
        10'd1011: TDATA = 39'b100010001001100010111000010110110100110;
        10'd1012: TDATA = 39'b100010001000011010111000000100100111010;
        10'd1013: TDATA = 39'b100010000111101010110111111000011110111;
        10'd1014: TDATA = 39'b100010000110100010110111100110010011011;
        10'd1015: TDATA = 39'b100010000101011010110111010100001001000;
        10'd1016: TDATA = 39'b100010000100010010110111000010000000000;
        10'd1017: TDATA = 39'b100010000011001010110110101111111000000;
        10'd1018: TDATA = 39'b100010000010000010110110011101110001010;
        10'd1019: TDATA = 39'b100010000000111010110110001011101011110;
        10'd1020: TDATA = 39'b100010000000001010110101111111101000110;
        10'd1021: TDATA = 39'b100001111111000010110101101101100101010;
        10'd1022: TDATA = 39'b100001111101111010110101011011100010111;
        10'd1023: TDATA = 39'b100001111100110010110101001001100001110;
	endcase
    end
    endfunction

    reg [7:0] ey_reg1,ey_reg2;
    reg [14:0] thalf_x0_reg;
    reg [22:0] mx_reg1,mx_reg2,mr_reg;
    reg [23:0] half_ax03_reg;

    // stage1
    wire odd_flag;
    wire [7:0] ex;
    wire [22:0] mx;
    wire [11:0] index;
    assign odd_flag = x[23];
    assign ex = x[30:23];
    assign mx = x[22:0];
    assign index = x[23:14];

    wire [38:0] tdata;
    assign tdata = TDATA(index);

    wire [14:0] thalf_x0;
    wire [23:0] half_x03;
    assign thalf_x0 = tdata[38:24];
    assign half_x03 = tdata[23:0];

    wire [7:0] ey;
    assign ey = (ex == 0) ? 0: (8'd63 + {1'b0,ex[7:1]} + odd_flag - (x[23:3] == {1'b1,20'b0} & x[2:0] < 3'd6));

    wire [47:0] half_ax03;
    assign half_ax03 = {1'b1,mx} * half_x03;

    // stage2
    wire [24:0] mra;
    assign mra = {thalf_x0_reg,10'b0} - {1'b0,half_ax03_reg};

    wire [22:0] mr;
    assign mr = mra[22:0];

    // stage 3
    wire [47:0] mya;
    assign mya = {1'b1,mr_reg} * {1'b1,mx_reg2};

    wire [22:0] my;
    assign my = (mya[47:47]) ? mya[46:24]: mya[45:23];

    assign y = {1'b0,ey_reg2,my};

    always @(posedge clk) begin
        // stage1
        ey_reg1 <= ey;
        mx_reg1 <= mx;
        thalf_x0_reg <= thalf_x0;
        half_ax03_reg <= half_ax03[47:24];
        // stage2
        ey_reg2 <= ey_reg1;
        mr_reg <= mr;
        mx_reg2 <= mx_reg1;
    end

    always @(negedge rstn) begin
        ey_reg1 <= 0;
        ey_reg2 <= 0;
        thalf_x0_reg <= 0;
        mx_reg1 <= 0;
        mx_reg2 <= 0;
        mr_reg <= 0;
        half_ax03_reg <= 0;
    end

endmodule
